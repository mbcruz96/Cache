
parameter SIZE = 20000;
module trace_addr(
    reg[31:0] test_addrs[0:SIZE-1]);
    
    assign test_addrs = 
    {
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034514,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034514,
    48'h00000400ed7b4,
    48'h00000400ed7b8,
    48'h000007b034400,
    48'h0000040020468,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfb0,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfb0,
    48'h00000400ed7c0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c18,
    48'h0000040045c18,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004002060c,
    48'h0000040020344,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b0344fc,
    48'h0000040020608,
    48'h000004002060c,
    48'h000004000e43c,
    48'h000007b0344fc,
    48'h000007b0344fc,
    48'h0000040059918,
    48'h000007b0337fc,
    48'h000007b0344fc,
    48'h00000400597c0,
    48'h0000040020608,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b034504,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b034504,
    48'h000007b0345b0,
    48'h000007b0345ac,
    48'h000007b0345a8,
    48'h000004002060c,
    48'h000004000e43c,
    48'h000007b0345b4,
    48'h000007b0345b4,
    48'h0000040059914,
    48'h00000400d602c,
    48'h000007b0345b0,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e5434,
    48'h00000400e5438,
    48'h000007b0345ac,
    48'h000007b0345cc,
    48'h000007b0345cc,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032344,
    48'h000007b0345a8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e53e4,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e5408,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b03463c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70c0,
    48'h000007b03464c,
    48'h000007b034648,
    48'h000007b034644,
    48'h000007b03464c,
    48'h000007b034648,
    48'h000007b034644,
    48'h000007b0337fc,
    48'h000007b03463c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bfc,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70bc,
    48'h00000400e70c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70d8,
    48'h00000400e70d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345b0,
    48'h00000400e53e0,
    48'h000007b0345a8,
    48'h000007b034400,
    48'h00000400ed790,
    48'h000007b034404,
    48'h00000400ed794,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004002078c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032348,
    48'h0000040020628,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h000004002079c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03438c,
    48'h000007b03438c,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h000007b03447c,
    48'h000004002078c,
    48'h0000040020610,
    48'h000007b0337fc,
    48'h0000040020614,
    48'h000004000e43c,
    48'h000007b03447c,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b034534,
    48'h0000040020610,
    48'h0000040020614,
    48'h000004000e43c,
    48'h000007b03453c,
    48'h000007b03453c,
    48'h0000040059918,
    48'h000007b0337fc,
    48'h0000040020610,
    48'h00000400e5434,
    48'h00000400e53e8,
    48'h000007b03453c,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b0345f8,
    48'h000007b0345f4,
    48'h000007b0345f0,
    48'h0000040020748,
    48'h000007b0345ec,
    48'h0000040058f58,
    48'h000007b0345ec,
    48'h000007b0345e8,
    48'h000007b034538,
    48'h00000400e5400,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf4,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6aac,
    48'h00000400e6ab4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6acc,
    48'h000007b034534,
    48'h00000400e6acc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034534,
    48'h00000400e5404,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf8,
    48'h00000400321e8,
    48'h0000040032328,
    48'h00000400e6db4,
    48'h00000400e6dbc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032328,
    48'h00000400e6dd4,
    48'h000007b0345f8,
    48'h00000400e6dd4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f8,
    48'h000007b0337fc,
    48'h00000400e5418,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bec,
    48'h00000400321e8,
    48'h000004003231c,
    48'h00000400e649c,
    48'h00000400e64a4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003231c,
    48'h00000400e64bc,
    48'h000007b0345fc,
    48'h00000400e64bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345fc,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b034694,
    48'h000007b034690,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h0000040059770,
    48'h000007b034698,
    48'h0000040059774,
    48'h000007b03469c,
    48'h0000040059778,
    48'h000007b0346a0,
    48'h000004005977c,
    48'h000007b0346a4,
    48'h0000040059780,
    48'h000007b0346a8,
    48'h0000040059784,
    48'h000007b0346ac,
    48'h0000040059788,
    48'h000007b0346b0,
    48'h000004005978c,
    48'h000007b0346b4,
    48'h0000040059790,
    48'h000007b0346b8,
    48'h0000040059794,
    48'h000007b0346bc,
    48'h00000400e5418,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003231c,
    48'h00000400e64a4,
    48'h000007b034694,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034694,
    48'h00000400e5418,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bec,
    48'h00000400321e8,
    48'h000004003231c,
    48'h00000400e649c,
    48'h00000400e64a4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003231c,
    48'h00000400e64bc,
    48'h000007b034690,
    48'h00000400e64bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b03477c,
    48'h000007b034778,
    48'h000007b034754,
    48'h000007b034750,
    48'h000007b0346a8,
    48'h000007b034690,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076190,
    48'h000007b034750,
    48'h0000040076190,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346b8,
    48'h000007b034750,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994a0,
    48'h000007b034778,
    48'h00000400994a0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034534,
    48'h000007b034778,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034804,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03480c,
    48'h000007b03480c,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h000007b034904,
    48'h0000040020054,
    48'h000007b034904,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034804,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h000007b034534,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h000007b034534,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000007b034534,
    48'h000004003bfb4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034804,
    48'h000007b034754,
    48'h000007b034804,
    48'h000007b034804,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000007b034534,
    48'h000004003234c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034778,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03483c,
    48'h000007b034754,
    48'h000007b0337fc,
    48'h000007b0346a8,
    48'h000007b034690,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076190,
    48'h000007b03483c,
    48'h0000040076190,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346b4,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034834,
    48'h000007b0337fc,
    48'h000007b034698,
    48'h000007b034754,
    48'h000007b034698,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034754,
    48'h00000400edc7c,
    48'h00000400edc80,
    48'h000007b034534,
    48'h0000040020468,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfb4,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfb4,
    48'h00000400edc88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c1c,
    48'h0000040045c1c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034778,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400e53f8,
    48'h00000400e53f4,
    48'h000007b0337fc,
    48'h00000400e5400,
    48'h000007b034534,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf4,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6aac,
    48'h00000400e6ab4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03473c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6acc,
    48'h00000400e6acc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400e5408,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70c0,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bfc,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70bc,
    48'h00000400e70c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70d8,
    48'h00000400e70d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400e5404,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf8,
    48'h00000400321e8,
    48'h0000040032328,
    48'h00000400e6db4,
    48'h00000400e6dbc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03473c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032328,
    48'h00000400e6dd4,
    48'h00000400e6dd4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400597c0,
    48'h00000400e53d4,
    48'h00000400e53c8,
    48'h00000400e5414,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c08,
    48'h00000400321e8,
    48'h0000040032338,
    48'h00000400ed254,
    48'h00000400ed25c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032338,
    48'h00000400ed274,
    48'h000007b03468c,
    48'h00000400ed274,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03468c,
    48'h000007b034534,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003234c,
    48'h000007b034688,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034534,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003234c,
    48'h00000400edc84,
    48'h000007b034684,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034688,
    48'h000007b034684,
    48'h00000400edc98,
    48'h000007b034684,
    48'h00000400edca0,
    48'h000007b034684,
    48'h00000400edca8,
    48'h000007b034684,
    48'h00000400edcb0,
    48'h000007b034684,
    48'h00000400edcb8,
    48'h000007b034684,
    48'h00000400edcc0,
    48'h000007b034684,
    48'h00000400edcc8,
    48'h000007b034684,
    48'h00000400edcd0,
    48'h000007b034684,
    48'h00000400edcd8,
    48'h000007b034684,
    48'h00000400edce0,
    48'h000007b034684,
    48'h00000400edce8,
    48'h000007b034684,
    48'h00000400edcf0,
    48'h000007b034684,
    48'h00000400edcf8,
    48'h000007b034684,
    48'h00000400edd00,
    48'h000007b034684,
    48'h00000400edd08,
    48'h000007b034684,
    48'h00000400edd10,
    48'h000007b034684,
    48'h00000400edd18,
    48'h000007b034684,
    48'h00000400edd20,
    48'h000007b034684,
    48'h00000400edd28,
    48'h000007b034684,
    48'h00000400edd30,
    48'h000007b034684,
    48'h00000400edd38,
    48'h000007b034684,
    48'h00000400edd40,
    48'h000007b034684,
    48'h00000400edd48,
    48'h000007b034684,
    48'h00000400edd50,
    48'h000007b034684,
    48'h00000400edd58,
    48'h000007b034684,
    48'h00000400edd60,
    48'h000007b034684,
    48'h00000400edd68,
    48'h000007b034684,
    48'h00000400edd70,
    48'h000007b034684,
    48'h00000400edd78,
    48'h000007b034684,
    48'h00000400edd80,
    48'h000007b034684,
    48'h00000400edd88,
    48'h000007b034684,
    48'h00000400edd90,
    48'h000007b034684,
    48'h00000400edd98,
    48'h000007b034684,
    48'h00000400edda0,
    48'h000007b034684,
    48'h00000400edda8,
    48'h000007b034684,
    48'h00000400eddb0,
    48'h000007b034684,
    48'h00000400eddb8,
    48'h000007b034684,
    48'h00000400eddc0,
    48'h000007b034684,
    48'h00000400eddc8,
    48'h000007b034684,
    48'h00000400eddd0,
    48'h000007b034684,
    48'h00000400eddd8,
    48'h000007b034684,
    48'h00000400edde0,
    48'h000007b034684,
    48'h00000400edde8,
    48'h000007b034684,
    48'h00000400eddf0,
    48'h000007b034684,
    48'h00000400eddf8,
    48'h000007b034684,
    48'h00000400ede00,
    48'h000007b034684,
    48'h00000400ede08,
    48'h000007b034684,
    48'h00000400ede10,
    48'h000007b034684,
    48'h00000400ede18,
    48'h000007b034684,
    48'h00000400ede20,
    48'h000007b034684,
    48'h00000400ede28,
    48'h000007b034684,
    48'h00000400ede30,
    48'h000007b034684,
    48'h00000400ede38,
    48'h000007b034684,
    48'h00000400ede40,
    48'h000007b034684,
    48'h00000400ede48,
    48'h000007b034684,
    48'h00000400ede50,
    48'h000007b034684,
    48'h00000400ede58,
    48'h000007b034684,
    48'h00000400ede60,
    48'h000007b034684,
    48'h00000400ede68,
    48'h000007b034684,
    48'h00000400ede70,
    48'h000007b034684,
    48'h00000400ede78,
    48'h000007b034684,
    48'h00000400ede80,
    48'h000007b034684,
    48'h00000400ede88,
    48'h000007b034684,
    48'h00000400ede90,
    48'h000007b034684,
    48'h00000400ede98,
    48'h000007b034684,
    48'h00000400edea0,
    48'h000007b034684,
    48'h00000400edea8,
    48'h000007b034684,
    48'h00000400edeb0,
    48'h000007b034684,
    48'h00000400edeb8,
    48'h000007b034684,
    48'h00000400edec0,
    48'h000007b034684,
    48'h00000400edec8,
    48'h000007b034684,
    48'h00000400eded0,
    48'h000007b034684,
    48'h00000400eded8,
    48'h000007b034684,
    48'h00000400edee0,
    48'h000007b034684,
    48'h00000400edee8,
    48'h000007b034684,
    48'h00000400edef0,
    48'h000007b034684,
    48'h00000400edef8,
    48'h000007b034684,
    48'h00000400edf00,
    48'h000007b034684,
    48'h00000400edf08,
    48'h000007b034684,
    48'h00000400edf10,
    48'h000007b034684,
    48'h00000400edf18,
    48'h000007b034684,
    48'h00000400edf20,
    48'h000007b034684,
    48'h00000400edf28,
    48'h000007b034684,
    48'h00000400edf30,
    48'h000007b034684,
    48'h00000400edf38,
    48'h000007b034684,
    48'h00000400edf40,
    48'h000007b034684,
    48'h00000400edf48,
    48'h000007b034684,
    48'h00000400edf50,
    48'h000007b034684,
    48'h00000400edf58,
    48'h000007b034684,
    48'h00000400edf60,
    48'h000007b034684,
    48'h00000400edf68,
    48'h000007b034684,
    48'h00000400edf70,
    48'h000007b034684,
    48'h00000400edf78,
    48'h000007b034684,
    48'h00000400edf80,
    48'h000007b034684,
    48'h00000400edf88,
    48'h000007b034684,
    48'h00000400edf90,
    48'h000007b034684,
    48'h00000400edf98,
    48'h000007b034684,
    48'h00000400edfa0,
    48'h000007b034684,
    48'h00000400edfa8,
    48'h000007b034684,
    48'h00000400edfb0,
    48'h000007b034684,
    48'h00000400edfb8,
    48'h000007b034684,
    48'h00000400edfc0,
    48'h000007b034684,
    48'h00000400edfc8,
    48'h000007b034684,
    48'h00000400edfd0,
    48'h000007b034684,
    48'h00000400edfd8,
    48'h000007b034684,
    48'h00000400edfe0,
    48'h000007b034684,
    48'h00000400edfe8,
    48'h000007b034684,
    48'h00000400edff0,
    48'h000007b034684,
    48'h00000400edff8,
    48'h000007b034684,
    48'h00000400ee000,
    48'h000007b034684,
    48'h00000400ee008,
    48'h000007b034684,
    48'h00000400ee010,
    48'h000007b034684,
    48'h00000400ee018,
    48'h000007b034684,
    48'h00000400ee020,
    48'h000007b034684,
    48'h00000400ee028,
    48'h000007b034684,
    48'h00000400ee030,
    48'h000007b034684,
    48'h00000400ee038,
    48'h000007b034684,
    48'h00000400ee040,
    48'h000007b034684,
    48'h00000400ee048,
    48'h000007b034684,
    48'h00000400ee050,
    48'h000007b034684,
    48'h00000400ee058,
    48'h000007b034684,
    48'h00000400ee060,
    48'h000007b034684,
    48'h00000400ee068,
    48'h000007b034684,
    48'h00000400ee070,
    48'h000007b034684,
    48'h00000400ee078,
    48'h000007b034684,
    48'h00000400ee080,
    48'h000007b034684,
    48'h00000400ee088,
    48'h000007b034684,
    48'h00000400ee090,
    48'h000007b034684,
    48'h00000400ee098,
    48'h000007b034684,
    48'h00000400ee0a0,
    48'h000007b034684,
    48'h00000400ee0a8,
    48'h000007b034684,
    48'h00000400ee0b0,
    48'h000007b034684,
    48'h00000400ee0b8,
    48'h000007b034684,
    48'h00000400ee0c0,
    48'h000007b034684,
    48'h00000400ee0c8,
    48'h000007b034684,
    48'h00000400ee0d0,
    48'h000007b034684,
    48'h00000400ee0d8,
    48'h000007b034684,
    48'h00000400ee0e0,
    48'h000007b034684,
    48'h00000400ee0e8,
    48'h000007b034684,
    48'h00000400ee0f0,
    48'h000007b034684,
    48'h00000400ee0f8,
    48'h000007b034684,
    48'h00000400ee100,
    48'h000007b034684,
    48'h00000400ee108,
    48'h000007b034684,
    48'h00000400ee110,
    48'h000007b034684,
    48'h00000400ee118,
    48'h000007b034684,
    48'h00000400ee120,
    48'h000007b034684,
    48'h00000400ee128,
    48'h000007b034684,
    48'h00000400ee130,
    48'h000007b034684,
    48'h00000400ee138,
    48'h000007b034684,
    48'h00000400ee140,
    48'h000007b034684,
    48'h00000400ee148,
    48'h000007b034684,
    48'h00000400ee150,
    48'h000007b034684,
    48'h00000400ee158,
    48'h000007b034684,
    48'h00000400ee160,
    48'h000007b034684,
    48'h00000400ee168,
    48'h000007b034684,
    48'h00000400ee170,
    48'h000007b034684,
    48'h00000400ee178,
    48'h000007b034684,
    48'h00000400ee180,
    48'h000007b034684,
    48'h00000400ee188,
    48'h000007b034684,
    48'h00000400ee190,
    48'h000007b034684,
    48'h00000400ee198,
    48'h000007b034684,
    48'h00000400ee1a0,
    48'h000007b034684,
    48'h00000400ee1a8,
    48'h000007b034684,
    48'h00000400ee1b0,
    48'h000007b034684,
    48'h00000400ee1b8,
    48'h000007b034684,
    48'h00000400ee1c0,
    48'h000007b034684,
    48'h00000400ee1c8,
    48'h000007b034684,
    48'h00000400ee1d0,
    48'h000007b034684,
    48'h00000400ee1d8,
    48'h000007b034684,
    48'h00000400ee1e0,
    48'h000007b034684,
    48'h00000400ee1e8,
    48'h000007b034684,
    48'h00000400ee1f0,
    48'h000007b034684,
    48'h00000400ee1f8,
    48'h000007b034684,
    48'h00000400ee200,
    48'h000007b034684,
    48'h00000400ee208,
    48'h000007b034684,
    48'h00000400ee210,
    48'h000007b034684,
    48'h00000400ee218,
    48'h000007b034684,
    48'h00000400ee220,
    48'h000007b034684,
    48'h00000400ee228,
    48'h000007b034684,
    48'h00000400ee230,
    48'h000007b034684,
    48'h00000400ee238,
    48'h000007b034684,
    48'h00000400ee240,
    48'h000007b034684,
    48'h00000400ee248,
    48'h000007b034684,
    48'h00000400ee250,
    48'h000007b034684,
    48'h00000400ee258,
    48'h000007b034684,
    48'h00000400ee260,
    48'h000007b034684,
    48'h00000400ee268,
    48'h000007b034684,
    48'h00000400ee270,
    48'h000007b034684,
    48'h00000400ee278,
    48'h000007b034684,
    48'h00000400ee280,
    48'h000007b034684,
    48'h00000400ee288,
    48'h000007b034684,
    48'h00000400ee290,
    48'h000007b034684,
    48'h00000400ee298,
    48'h000007b034684,
    48'h00000400ee2a0,
    48'h000007b034684,
    48'h00000400ee2a8,
    48'h000007b034684,
    48'h00000400ee2b0,
    48'h000007b034684,
    48'h00000400ee2b8,
    48'h000007b034684,
    48'h00000400ee2c0,
    48'h000007b034684,
    48'h00000400ee2c8,
    48'h000007b034684,
    48'h00000400ee2d0,
    48'h000007b034684,
    48'h00000400ee2d8,
    48'h000007b034684,
    48'h00000400ee2e0,
    48'h000007b034684,
    48'h00000400ee2e8,
    48'h000007b034684,
    48'h00000400ee2f0,
    48'h000007b034684,
    48'h00000400ee2f8,
    48'h000007b034684,
    48'h00000400ee300,
    48'h000007b034684,
    48'h00000400ee308,
    48'h000007b034684,
    48'h00000400ee310,
    48'h000007b034684,
    48'h00000400ee318,
    48'h000007b034684,
    48'h00000400ee320,
    48'h000007b034684,
    48'h00000400ee328,
    48'h000007b034684,
    48'h00000400ee330,
    48'h000007b034684,
    48'h00000400ee338,
    48'h000007b034684,
    48'h00000400ee340,
    48'h000007b034684,
    48'h00000400ee348,
    48'h000007b034684,
    48'h00000400ee350,
    48'h000007b034684,
    48'h00000400ee358,
    48'h000007b034684,
    48'h00000400ee360,
    48'h000007b034684,
    48'h00000400ee368,
    48'h000007b034684,
    48'h00000400ee370,
    48'h000007b034684,
    48'h00000400ee378,
    48'h000007b034684,
    48'h00000400ee380,
    48'h000007b034684,
    48'h00000400ee388,
    48'h000007b034684,
    48'h00000400ee390,
    48'h000007b034684,
    48'h00000400ee398,
    48'h000007b034684,
    48'h00000400ee3a0,
    48'h000007b034684,
    48'h00000400ee3a8,
    48'h000007b034684,
    48'h00000400ee3b0,
    48'h000007b034684,
    48'h00000400ee3b8,
    48'h000007b034684,
    48'h00000400ee3c0,
    48'h000007b034684,
    48'h00000400ee3c8,
    48'h000007b034684,
    48'h00000400ee3d0,
    48'h000007b034684,
    48'h00000400ee3d8,
    48'h000007b034684,
    48'h00000400ee3e0,
    48'h000007b034684,
    48'h00000400ee3e8,
    48'h000007b034684,
    48'h00000400ee3f0,
    48'h000007b034684,
    48'h00000400ee3f8,
    48'h000007b034684,
    48'h00000400ee400,
    48'h000007b034684,
    48'h00000400ee408,
    48'h000007b034684,
    48'h00000400ee410,
    48'h000007b034684,
    48'h00000400ee418,
    48'h000007b034684,
    48'h00000400ee420,
    48'h000007b034684,
    48'h00000400ee428,
    48'h000007b034684,
    48'h00000400ee430,
    48'h000007b034684,
    48'h00000400ee438,
    48'h000007b034684,
    48'h00000400ee440,
    48'h000007b034684,
    48'h00000400ee448,
    48'h000007b034684,
    48'h00000400ee450,
    48'h000007b034684,
    48'h00000400ee458,
    48'h000007b034684,
    48'h00000400ee460,
    48'h000007b034684,
    48'h00000400ee468,
    48'h000007b034684,
    48'h00000400ee470,
    48'h000007b034684,
    48'h00000400ee478,
    48'h000007b034684,
    48'h00000400ee480,
    48'h000007b034684,
    48'h00000400ee488,
    48'h000007b034684,
    48'h00000400ee490,
    48'h000007b034684,
    48'h00000400ee498,
    48'h000007b034684,
    48'h00000400ee4a0,
    48'h000007b034684,
    48'h00000400ee4a8,
    48'h000007b034684,
    48'h00000400ee4b0,
    48'h000007b034684,
    48'h00000400ee4b8,
    48'h000007b034684,
    48'h00000400ee4c0,
    48'h000007b034684,
    48'h00000400ee4c8,
    48'h000007b034684,
    48'h00000400ee4d0,
    48'h000007b034684,
    48'h00000400ee4d8,
    48'h000007b034684,
    48'h00000400ee4e0,
    48'h000007b034684,
    48'h00000400ee4e8,
    48'h000007b034684,
    48'h00000400ee4f0,
    48'h000007b034684,
    48'h00000400ee4f8,
    48'h000007b034684,
    48'h00000400ee500,
    48'h000007b034684,
    48'h00000400ee508,
    48'h000007b034684,
    48'h00000400ee510,
    48'h000007b034684,
    48'h00000400ee518,
    48'h000007b034684,
    48'h00000400ee520,
    48'h000007b034684,
    48'h00000400ee528,
    48'h000007b034684,
    48'h00000400ee530,
    48'h000007b034684,
    48'h00000400ee538,
    48'h000007b034684,
    48'h00000400ee540,
    48'h000007b034684,
    48'h00000400ee548,
    48'h000007b034684,
    48'h00000400ee550,
    48'h000007b034684,
    48'h00000400ee558,
    48'h000007b034684,
    48'h00000400ee560,
    48'h000007b034684,
    48'h00000400ee568,
    48'h000007b034684,
    48'h00000400ee570,
    48'h000007b034684,
    48'h00000400ee578,
    48'h000007b034684,
    48'h00000400ee580,
    48'h000007b034684,
    48'h00000400ee588,
    48'h000007b034684,
    48'h00000400ee590,
    48'h000007b034684,
    48'h00000400ee598,
    48'h000007b034684,
    48'h00000400ee5a0,
    48'h000007b034684,
    48'h00000400ee5a8,
    48'h000007b034684,
    48'h00000400ee5b0,
    48'h000007b034684,
    48'h00000400ee5b8,
    48'h000007b034684,
    48'h00000400ee5c0,
    48'h000007b034684,
    48'h00000400ee5c8,
    48'h000007b034684,
    48'h00000400ee5d0,
    48'h000007b034684,
    48'h00000400ee5d8,
    48'h000007b034684,
    48'h00000400ee5e0,
    48'h000007b034684,
    48'h00000400ee5e8,
    48'h000007b034684,
    48'h00000400ee5f0,
    48'h000007b034684,
    48'h00000400ee5f8,
    48'h000007b034684,
    48'h00000400ee600,
    48'h000007b034684,
    48'h00000400ee608,
    48'h000007b034684,
    48'h00000400ee610,
    48'h000007b034684,
    48'h00000400ee618,
    48'h000007b034684,
    48'h00000400ee620,
    48'h000007b034684,
    48'h00000400ee628,
    48'h000007b034684,
    48'h00000400ee630,
    48'h000007b034684,
    48'h00000400ee638,
    48'h000007b034684,
    48'h00000400ee640,
    48'h000007b034684,
    48'h00000400ee648,
    48'h000007b034684,
    48'h00000400ee650,
    48'h000007b034684,
    48'h00000400ee658,
    48'h000007b034684,
    48'h00000400ee660,
    48'h000007b034684,
    48'h00000400ee668,
    48'h000007b034684,
    48'h00000400ee670,
    48'h000007b034684,
    48'h00000400ee678,
    48'h000007b034684,
    48'h00000400ee680,
    48'h000007b034684,
    48'h00000400ee688,
    48'h000007b034684,
    48'h00000400ee690,
    48'h000007b034684,
    48'h00000400ee698,
    48'h000007b034684,
    48'h00000400ee6a0,
    48'h000007b034684,
    48'h00000400ee6a8,
    48'h000007b034684,
    48'h00000400ee6b0,
    48'h000007b034684,
    48'h00000400ee6b8,
    48'h000007b034684,
    48'h00000400ee6c0,
    48'h000007b034684,
    48'h00000400ee6c8,
    48'h000007b034684,
    48'h00000400ee6d0,
    48'h000007b034684,
    48'h00000400ee6d8,
    48'h000007b034684,
    48'h00000400ee6e0,
    48'h000007b034684,
    48'h00000400ee6e8,
    48'h000007b034684,
    48'h00000400ee6f0,
    48'h000007b034684,
    48'h00000400ee6f8,
    48'h000007b034684,
    48'h00000400ee700,
    48'h000007b034684,
    48'h00000400ee708,
    48'h000007b034684,
    48'h00000400ee710,
    48'h000007b034684,
    48'h00000400ee718,
    48'h000007b034684,
    48'h00000400ee720,
    48'h000007b034684,
    48'h00000400ee728,
    48'h000007b034684,
    48'h00000400ee730,
    48'h000007b034684,
    48'h00000400ee738,
    48'h000007b034684,
    48'h00000400ee740,
    48'h000007b034684,
    48'h00000400ee748,
    48'h000007b034684,
    48'h00000400ee750,
    48'h000007b034684,
    48'h00000400ee758,
    48'h000007b034684,
    48'h00000400ee760,
    48'h000007b034684,
    48'h00000400ee768,
    48'h000007b034684,
    48'h00000400ee770,
    48'h000007b034684,
    48'h00000400ee778,
    48'h000007b034684,
    48'h00000400ee780,
    48'h000007b034684,
    48'h00000400ee788,
    48'h000007b034684,
    48'h00000400ee790,
    48'h000007b034684,
    48'h00000400ee798,
    48'h000007b034684,
    48'h00000400ee7a0,
    48'h000007b034684,
    48'h00000400ee7a8,
    48'h000007b034684,
    48'h00000400ee7b0,
    48'h000007b034684,
    48'h00000400ee7b8,
    48'h000007b034684,
    48'h00000400ee7c0,
    48'h000007b034684,
    48'h00000400ee7c8,
    48'h000007b034684,
    48'h00000400ee7d0,
    48'h000007b034684,
    48'h00000400ee7d8,
    48'h000007b034684,
    48'h00000400ee7e0,
    48'h000007b034684,
    48'h00000400ee7e8,
    48'h000007b034684,
    48'h00000400ee7f0,
    48'h000007b034684,
    48'h00000400ee7f8,
    48'h000007b034684,
    48'h00000400ee800,
    48'h000007b034684,
    48'h00000400ee808,
    48'h000007b034684,
    48'h00000400ee810,
    48'h000007b034684,
    48'h00000400ee818,
    48'h000007b034684,
    48'h00000400ee820,
    48'h000007b034684,
    48'h00000400ee828,
    48'h000007b034684,
    48'h00000400ee830,
    48'h000007b034684,
    48'h00000400ee838,
    48'h000007b034684,
    48'h00000400ee840,
    48'h000007b034684,
    48'h00000400ee848,
    48'h000007b034684,
    48'h00000400ee850,
    48'h000007b034684,
    48'h00000400ee858,
    48'h000007b034684,
    48'h00000400ee860,
    48'h000007b034684,
    48'h00000400ee868,
    48'h000007b034684,
    48'h00000400ee870,
    48'h000007b034684,
    48'h00000400ee878,
    48'h000007b034684,
    48'h00000400ee880,
    48'h000007b034684,
    48'h00000400ee888,
    48'h000007b034684,
    48'h00000400ee890,
    48'h000007b034684,
    48'h00000400ee898,
    48'h000007b034684,
    48'h00000400ee8a0,
    48'h000007b034684,
    48'h00000400ee8a8,
    48'h000007b034684,
    48'h00000400ee8b0,
    48'h000007b034684,
    48'h00000400ee8b8,
    48'h000007b034684,
    48'h00000400ee8c0,
    48'h000007b034684,
    48'h00000400ee8c8,
    48'h000007b034684,
    48'h00000400ee8d0,
    48'h000007b034684,
    48'h00000400ee8d8,
    48'h000007b034684,
    48'h00000400ee8e0,
    48'h000007b034684,
    48'h00000400ee8e8,
    48'h000007b034684,
    48'h00000400ee8f0,
    48'h000007b034684,
    48'h00000400ee8f8,
    48'h000007b034684,
    48'h00000400ee900,
    48'h000007b034684,
    48'h00000400ee908,
    48'h000007b034684,
    48'h00000400ee910,
    48'h000007b034684,
    48'h00000400ee918,
    48'h000007b034684,
    48'h00000400ee920,
    48'h000007b034684,
    48'h00000400ee928,
    48'h000007b034684,
    48'h00000400ee930,
    48'h000007b034684,
    48'h00000400ee938,
    48'h000007b034684,
    48'h00000400ee940,
    48'h000007b034684,
    48'h00000400ee948,
    48'h000007b034684,
    48'h00000400ee950,
    48'h000007b034684,
    48'h00000400ee958,
    48'h000007b034684,
    48'h00000400ee960,
    48'h000007b034684,
    48'h00000400ee968,
    48'h000007b034684,
    48'h00000400ee970,
    48'h000007b034684,
    48'h00000400ee978,
    48'h000007b034684,
    48'h00000400ee980,
    48'h000007b034684,
    48'h00000400ee988,
    48'h000007b034684,
    48'h00000400ee990,
    48'h000007b034684,
    48'h00000400ee998,
    48'h000007b034684,
    48'h00000400ee9a0,
    48'h000007b034684,
    48'h00000400ee9a8,
    48'h000007b034684,
    48'h00000400ee9b0,
    48'h000007b034684,
    48'h00000400ee9b8,
    48'h000007b034684,
    48'h00000400ee9c0,
    48'h000007b034684,
    48'h00000400ee9c8,
    48'h000007b034684,
    48'h00000400ee9d0,
    48'h000007b034684,
    48'h00000400ee9d8,
    48'h000007b034684,
    48'h00000400ee9e0,
    48'h000007b034684,
    48'h00000400ee9e8,
    48'h000007b034684,
    48'h00000400ee9f0,
    48'h000007b034684,
    48'h00000400ee9f8,
    48'h000007b034684,
    48'h00000400eea00,
    48'h000007b034684,
    48'h00000400eea08,
    48'h000007b034684,
    48'h00000400eea10,
    48'h000007b034684,
    48'h00000400eea18,
    48'h000007b034684,
    48'h00000400eea20,
    48'h000007b034684,
    48'h00000400eea28,
    48'h000007b034684,
    48'h00000400eea30,
    48'h000007b034684,
    48'h00000400eea38,
    48'h000007b034684,
    48'h00000400eea40,
    48'h000007b034684,
    48'h00000400eea48,
    48'h000007b034684,
    48'h00000400eea50,
    48'h000007b034684,
    48'h00000400eea58,
    48'h000007b034684,
    48'h00000400eea60,
    48'h000007b034684,
    48'h00000400eea68,
    48'h000007b034684,
    48'h00000400eea70,
    48'h000007b034684,
    48'h00000400eea78,
    48'h000007b034684,
    48'h00000400eea80,
    48'h000007b034684,
    48'h00000400eea88,
    48'h000007b034684,
    48'h00000400eea90,
    48'h000007b034684,
    48'h00000400eea98,
    48'h000007b034684,
    48'h00000400eeaa0,
    48'h000007b034684,
    48'h00000400eeaa8,
    48'h000007b034684,
    48'h00000400eeab0,
    48'h000007b034684,
    48'h00000400eeab8,
    48'h000007b034684,
    48'h00000400eeac0,
    48'h000007b034684,
    48'h00000400eeac8,
    48'h000007b034684,
    48'h00000400eead0,
    48'h000007b034684,
    48'h00000400eead8,
    48'h000007b034684,
    48'h00000400eeae0,
    48'h000007b034684,
    48'h00000400eeae8,
    48'h000007b034684,
    48'h00000400eeaf0,
    48'h000007b034684,
    48'h00000400eeaf8,
    48'h000007b034684,
    48'h00000400eeb00,
    48'h000007b034684,
    48'h00000400eeb08,
    48'h000007b034684,
    48'h00000400eeb10,
    48'h000007b034684,
    48'h00000400eeb18,
    48'h000007b034684,
    48'h00000400eeb20,
    48'h000007b034684,
    48'h00000400eeb28,
    48'h000007b034684,
    48'h00000400eeb30,
    48'h000007b034684,
    48'h00000400eeb38,
    48'h000007b034684,
    48'h00000400eeb40,
    48'h000007b034684,
    48'h00000400eeb48,
    48'h000007b034684,
    48'h00000400eeb50,
    48'h000007b034684,
    48'h00000400eeb58,
    48'h000007b034684,
    48'h00000400eeb60,
    48'h000007b034684,
    48'h00000400eeb68,
    48'h000007b034684,
    48'h00000400eeb70,
    48'h000007b034684,
    48'h00000400eeb78,
    48'h000007b034684,
    48'h00000400eeb80,
    48'h000007b034684,
    48'h00000400eeb88,
    48'h000007b034684,
    48'h00000400eeb90,
    48'h000007b034684,
    48'h00000400eeb98,
    48'h000007b034684,
    48'h00000400eeba0,
    48'h000007b034684,
    48'h00000400eeba8,
    48'h000007b034684,
    48'h00000400eebb0,
    48'h000007b034684,
    48'h00000400eebb8,
    48'h000007b034684,
    48'h00000400eebc0,
    48'h000007b034684,
    48'h00000400eebc8,
    48'h000007b034684,
    48'h00000400eebd0,
    48'h000007b034684,
    48'h00000400eebd8,
    48'h000007b034684,
    48'h00000400eebe0,
    48'h000007b034684,
    48'h00000400eebe8,
    48'h000007b034684,
    48'h00000400eebf0,
    48'h000007b034684,
    48'h00000400eebf8,
    48'h000007b034684,
    48'h00000400eec00,
    48'h000007b034684,
    48'h00000400eec08,
    48'h000007b034684,
    48'h00000400eec10,
    48'h000007b034684,
    48'h00000400eec18,
    48'h000007b034684,
    48'h00000400eec20,
    48'h000007b034684,
    48'h00000400eec28,
    48'h000007b034684,
    48'h00000400eec30,
    48'h000007b034684,
    48'h00000400eec38,
    48'h000007b034684,
    48'h00000400eec40,
    48'h000007b034684,
    48'h00000400eec48,
    48'h000007b034684,
    48'h00000400eec50,
    48'h000007b034684,
    48'h00000400eec58,
    48'h000007b034684,
    48'h00000400eec60,
    48'h000007b034684,
    48'h00000400eec68,
    48'h000007b034684,
    48'h00000400eec70,
    48'h000007b034684,
    48'h00000400eec78,
    48'h000007b034684,
    48'h00000400eec80,
    48'h000007b034684,
    48'h00000400eec88,
    48'h000007b034684,
    48'h00000400eec90,
    48'h000007b034684,
    48'h00000400eec98,
    48'h000007b034684,
    48'h00000400eeca0,
    48'h000007b034684,
    48'h00000400eeca8,
    48'h000007b034684,
    48'h00000400eecb0,
    48'h000007b034684,
    48'h00000400eecb8,
    48'h000007b034684,
    48'h00000400eecc0,
    48'h000007b034684,
    48'h00000400eecc8,
    48'h000007b034684,
    48'h00000400eecd0,
    48'h000007b034684,
    48'h00000400eecd8,
    48'h000007b034684,
    48'h00000400eece0,
    48'h000007b034684,
    48'h00000400eece8,
    48'h000007b034684,
    48'h00000400eecf0,
    48'h000007b034684,
    48'h00000400eecf8,
    48'h000007b034684,
    48'h00000400eed00,
    48'h000007b034684,
    48'h00000400eed08,
    48'h000007b034684,
    48'h00000400eed10,
    48'h000007b034684,
    48'h00000400eed18,
    48'h000007b034684,
    48'h00000400eed20,
    48'h000007b034684,
    48'h00000400eed28,
    48'h000007b034684,
    48'h00000400eed30,
    48'h000007b034684,
    48'h00000400eed38,
    48'h000007b034684,
    48'h00000400eed40,
    48'h000007b034684,
    48'h00000400eed48,
    48'h000007b034684,
    48'h00000400eed50,
    48'h000007b034684,
    48'h00000400eed58,
    48'h000007b034684,
    48'h00000400eed60,
    48'h000007b034684,
    48'h00000400eed68,
    48'h000007b034684,
    48'h00000400eed70,
    48'h000007b034684,
    48'h00000400eed78,
    48'h000007b034684,
    48'h00000400eed80,
    48'h000007b034684,
    48'h00000400eed88,
    48'h000007b034684,
    48'h00000400eed90,
    48'h000007b034684,
    48'h00000400eed98,
    48'h000007b034684,
    48'h00000400eeda0,
    48'h000007b034684,
    48'h00000400eeda8,
    48'h000007b034684,
    48'h00000400eedb0,
    48'h000007b034684,
    48'h00000400eedb8,
    48'h000007b034684,
    48'h00000400eedc0,
    48'h000007b034684,
    48'h00000400eedc8,
    48'h000007b034684,
    48'h00000400eedd0,
    48'h000007b034684,
    48'h00000400eedd8,
    48'h000007b034684,
    48'h00000400eede0,
    48'h000007b034684,
    48'h00000400eede8,
    48'h000007b034684,
    48'h00000400eedf0,
    48'h000007b034684,
    48'h00000400eedf8,
    48'h000007b034684,
    48'h00000400eee00,
    48'h000007b034684,
    48'h00000400eee08,
    48'h000007b034684,
    48'h00000400eee10,
    48'h000007b034684,
    48'h00000400eee18,
    48'h000007b034684,
    48'h00000400eee20,
    48'h000007b034684,
    48'h00000400eee28,
    48'h000007b034684,
    48'h00000400eee30,
    48'h000007b034684,
    48'h00000400eee38,
    48'h000007b034684,
    48'h00000400eee40,
    48'h000007b034684,
    48'h00000400eee48,
    48'h000007b034684,
    48'h00000400eee50,
    48'h000007b034684,
    48'h00000400eee58,
    48'h000007b034684,
    48'h00000400eee60,
    48'h000007b034684,
    48'h00000400eee68,
    48'h000007b034684,
    48'h00000400eee70,
    48'h000007b034684,
    48'h00000400eee78,
    48'h000007b034684,
    48'h00000400eee80,
    48'h000007b034684,
    48'h00000400eee88,
    48'h000007b034684,
    48'h00000400eee90,
    48'h000007b034684,
    48'h00000400eee98,
    48'h000007b034684,
    48'h00000400eeea0,
    48'h000007b034684,
    48'h00000400eeea8,
    48'h000007b034684,
    48'h00000400eeeb0,
    48'h000007b034684,
    48'h00000400eeeb8,
    48'h000007b034684,
    48'h00000400eeec0,
    48'h000007b034684,
    48'h00000400eeec8,
    48'h000007b034684,
    48'h00000400eeed0,
    48'h000007b034684,
    48'h00000400eeed8,
    48'h000007b034684,
    48'h00000400eeee0,
    48'h000007b034684,
    48'h00000400eeee8,
    48'h000007b034684,
    48'h00000400eeef0,
    48'h000007b034684,
    48'h00000400eeef8,
    48'h000007b034684,
    48'h00000400eef00,
    48'h000007b034684,
    48'h00000400eef08,
    48'h000007b034684,
    48'h00000400eef10,
    48'h000007b034684,
    48'h00000400eef18,
    48'h000007b034684,
    48'h00000400eef20,
    48'h000007b034684,
    48'h00000400eef28,
    48'h000007b034684,
    48'h00000400eef30,
    48'h000007b034684,
    48'h00000400eef38,
    48'h000007b034684,
    48'h00000400eef40,
    48'h000007b034684,
    48'h00000400eef48,
    48'h000007b034684,
    48'h00000400eef50,
    48'h000007b034684,
    48'h00000400eef58,
    48'h000007b034684,
    48'h00000400eef60,
    48'h000007b034684,
    48'h00000400eef68,
    48'h000007b034684,
    48'h00000400eef70,
    48'h000007b034684,
    48'h00000400eef78,
    48'h000007b034684,
    48'h00000400eef80,
    48'h000007b034684,
    48'h00000400eef88,
    48'h000007b034684,
    48'h00000400eef90,
    48'h000007b034684,
    48'h00000400eef98,
    48'h000007b034684,
    48'h00000400eefa0,
    48'h000007b034684,
    48'h00000400eefa8,
    48'h000007b034684,
    48'h00000400eefb0,
    48'h000007b034684,
    48'h00000400eefb8,
    48'h000007b034684,
    48'h00000400eefc0,
    48'h000007b034684,
    48'h00000400eefc8,
    48'h000007b034684,
    48'h00000400eefd0,
    48'h000007b034684,
    48'h00000400eefd8,
    48'h000007b034684,
    48'h00000400eefe0,
    48'h000007b034684,
    48'h00000400eefe8,
    48'h000007b034684,
    48'h00000400eeff0,
    48'h000007b034684,
    48'h00000400eeff8,
    48'h000007b034684,
    48'h00000400ef000,
    48'h000007b034684,
    48'h00000400ef008,
    48'h000007b034684,
    48'h00000400ef010,
    48'h000007b034684,
    48'h00000400ef018,
    48'h000007b034684,
    48'h00000400ef020,
    48'h000007b034684,
    48'h00000400ef028,
    48'h000007b034684,
    48'h00000400ef030,
    48'h000007b034684,
    48'h00000400ef038,
    48'h000007b034684,
    48'h00000400ef040,
    48'h000007b034684,
    48'h00000400ef048,
    48'h000007b034684,
    48'h00000400ef050,
    48'h000007b034684,
    48'h00000400ef058,
    48'h000007b034684,
    48'h00000400ef060,
    48'h000007b034684,
    48'h00000400ef068,
    48'h000007b034684,
    48'h00000400ef070,
    48'h000007b034684,
    48'h00000400ef078,
    48'h000007b034684,
    48'h00000400ef080,
    48'h000007b034684,
    48'h00000400ef088,
    48'h000007b034684,
    48'h00000400ef090,
    48'h000007b034684,
    48'h00000400ef098,
    48'h000007b034684,
    48'h00000400ef0a0,
    48'h000007b034684,
    48'h00000400ef0a8,
    48'h000007b034684,
    48'h00000400ef0b0,
    48'h000007b034684,
    48'h00000400ef0b8,
    48'h000007b034684,
    48'h00000400ef0c0,
    48'h000007b034684,
    48'h00000400ef0c8,
    48'h000007b034684,
    48'h00000400ef0d0,
    48'h000007b034684,
    48'h00000400ef0d8,
    48'h000007b034684,
    48'h00000400ef0e0,
    48'h000007b034684,
    48'h00000400ef0e8,
    48'h000007b034684,
    48'h00000400ef0f0,
    48'h000007b034684,
    48'h00000400ef0f8,
    48'h000007b034684,
    48'h00000400ef100,
    48'h000007b034684,
    48'h00000400ef108,
    48'h000007b034684,
    48'h00000400ef110,
    48'h000007b034684,
    48'h00000400ef118,
    48'h000007b034684,
    48'h00000400ef120,
    48'h000007b034684,
    48'h00000400ef128,
    48'h000007b034684,
    48'h00000400ef130,
    48'h000007b034684,
    48'h00000400ef138,
    48'h000007b034684,
    48'h00000400ef140,
    48'h000007b034684,
    48'h00000400ef148,
    48'h000007b034684,
    48'h00000400ef150,
    48'h000007b034684,
    48'h00000400ef158,
    48'h000007b034684,
    48'h00000400ef160,
    48'h000007b034684,
    48'h00000400ef168,
    48'h000007b034684,
    48'h00000400ef170,
    48'h000007b034684,
    48'h00000400ef178,
    48'h000007b034684,
    48'h00000400ef180,
    48'h000007b034684,
    48'h00000400ef188,
    48'h000007b034684,
    48'h00000400ef190,
    48'h000007b034684,
    48'h00000400ef198,
    48'h000007b034684,
    48'h00000400ef1a0,
    48'h000007b034684,
    48'h00000400ef1a8,
    48'h000007b034684,
    48'h00000400ef1b0,
    48'h000007b034684,
    48'h00000400ef1b8,
    48'h000007b034684,
    48'h00000400ef1c0,
    48'h000007b034684,
    48'h00000400ef1c8,
    48'h000007b034684,
    48'h00000400ef1d0,
    48'h000007b034684,
    48'h00000400ef1d8,
    48'h000007b034684,
    48'h00000400ef1e0,
    48'h000007b034684,
    48'h00000400ef1e8,
    48'h000007b034684,
    48'h00000400ef1f0,
    48'h000007b034684,
    48'h00000400ef1f8,
    48'h000007b034684,
    48'h00000400ef200,
    48'h000007b034684,
    48'h00000400ef208,
    48'h000007b034684,
    48'h00000400ef210,
    48'h000007b034684,
    48'h00000400ef218,
    48'h000007b034684,
    48'h00000400ef220,
    48'h000007b034684,
    48'h00000400ef228,
    48'h000007b034684,
    48'h00000400ef230,
    48'h000007b034684,
    48'h00000400ef238,
    48'h000007b034684,
    48'h00000400ef240,
    48'h000007b034684,
    48'h00000400ef248,
    48'h000007b034684,
    48'h00000400ef250,
    48'h000007b034684,
    48'h00000400ef258,
    48'h000007b034684,
    48'h00000400ef260,
    48'h000007b034684,
    48'h00000400ef268,
    48'h000007b034684,
    48'h00000400ef270,
    48'h000007b034684,
    48'h00000400ef278,
    48'h000007b034684,
    48'h00000400ef280,
    48'h000007b034684,
    48'h00000400ef288,
    48'h000007b034684,
    48'h00000400ef290,
    48'h000007b034684,
    48'h00000400ef298,
    48'h000007b034684,
    48'h00000400ef2a0,
    48'h000007b034684,
    48'h00000400ef2a8,
    48'h000007b034684,
    48'h00000400ef2b0,
    48'h000007b034684,
    48'h00000400ef2b8,
    48'h000007b034684,
    48'h00000400ef2c0,
    48'h000007b034684,
    48'h00000400ef2c8,
    48'h000007b034684,
    48'h00000400ef2d0,
    48'h000007b034684,
    48'h00000400ef2d8,
    48'h000007b034684,
    48'h00000400ef2e0,
    48'h000007b034684,
    48'h00000400ef2e8,
    48'h000007b034684,
    48'h00000400ef2f0,
    48'h000007b034684,
    48'h00000400ef2f8,
    48'h000007b034684,
    48'h00000400ef300,
    48'h000007b034684,
    48'h00000400ef308,
    48'h000007b034684,
    48'h00000400ef310,
    48'h000007b034684,
    48'h00000400ef318,
    48'h000007b034684,
    48'h00000400ef320,
    48'h000007b034684,
    48'h00000400ef328,
    48'h000007b034684,
    48'h00000400ef330,
    48'h000007b034684,
    48'h00000400ef338,
    48'h000007b034684,
    48'h00000400ef340,
    48'h000007b034684,
    48'h00000400ef348,
    48'h000007b034684,
    48'h00000400ef350,
    48'h000007b034684,
    48'h00000400ef358,
    48'h000007b034684,
    48'h00000400ef360,
    48'h000007b034684,
    48'h00000400ef368,
    48'h000007b034684,
    48'h00000400ef370,
    48'h000007b034684,
    48'h00000400ef378,
    48'h000007b034684,
    48'h00000400ef380,
    48'h000007b034684,
    48'h00000400ef388,
    48'h000007b034684,
    48'h00000400ef390,
    48'h000007b034684,
    48'h00000400ef398,
    48'h000007b034684,
    48'h00000400ef3a0,
    48'h000007b034684,
    48'h00000400ef3a8,
    48'h000007b034684,
    48'h00000400ef3b0,
    48'h000007b034684,
    48'h00000400ef3b8,
    48'h000007b034684,
    48'h00000400ef3c0,
    48'h000007b034684,
    48'h00000400ef3c8,
    48'h000007b034684,
    48'h00000400ef3d0,
    48'h000007b034684,
    48'h00000400ef3d8,
    48'h000007b034684,
    48'h00000400ef3e0,
    48'h000007b034684,
    48'h00000400ef3e8,
    48'h000007b034684,
    48'h00000400ef3f0,
    48'h000007b034684,
    48'h00000400ef3f8,
    48'h000007b034684,
    48'h00000400ef400,
    48'h000007b034684,
    48'h00000400ef408,
    48'h000007b034684,
    48'h00000400ef410,
    48'h000007b034684,
    48'h00000400ef418,
    48'h000007b034684,
    48'h00000400ef420,
    48'h000007b034684,
    48'h00000400ef428,
    48'h000007b034684,
    48'h00000400ef430,
    48'h000007b034684,
    48'h00000400ef438,
    48'h000007b034684,
    48'h00000400ef440,
    48'h000007b034684,
    48'h00000400ef448,
    48'h000007b034684,
    48'h00000400ef450,
    48'h000007b034684,
    48'h00000400ef458,
    48'h000007b034684,
    48'h00000400ef460,
    48'h000007b034684,
    48'h00000400ef468,
    48'h000007b034684,
    48'h00000400ef470,
    48'h000007b034684,
    48'h00000400ef478,
    48'h000007b034684,
    48'h00000400ef480,
    48'h000007b034684,
    48'h00000400ef488,
    48'h000007b034684,
    48'h00000400ef490,
    48'h000007b034684,
    48'h00000400ef498,
    48'h000007b034684,
    48'h00000400ef4a0,
    48'h000007b034684,
    48'h00000400ef4a8,
    48'h000007b034684,
    48'h00000400ef4b0,
    48'h000007b034684,
    48'h00000400ef4b8,
    48'h000007b034684,
    48'h00000400ef4c0,
    48'h000007b034684,
    48'h00000400ef4c8,
    48'h000007b034684,
    48'h00000400ef4d0,
    48'h000007b034684,
    48'h00000400ef4d8,
    48'h000007b034684,
    48'h00000400ef4e0,
    48'h000007b034684,
    48'h00000400ef4e8,
    48'h000007b034684,
    48'h00000400ef4f0,
    48'h000007b034684,
    48'h00000400ef4f8,
    48'h000007b034684,
    48'h00000400ef500,
    48'h000007b034684,
    48'h00000400ef508,
    48'h000007b034684,
    48'h00000400ef510,
    48'h000007b034684,
    48'h00000400ef518,
    48'h000007b034684,
    48'h00000400ef520,
    48'h000007b034684,
    48'h00000400ef528,
    48'h000007b034684,
    48'h00000400ef530,
    48'h000007b034684,
    48'h00000400ef538,
    48'h000007b034684,
    48'h00000400ef540,
    48'h000007b034684,
    48'h00000400ef548,
    48'h000007b034684,
    48'h00000400ef550,
    48'h000007b034684,
    48'h00000400ef558,
    48'h000007b034684,
    48'h00000400ef560,
    48'h000007b034684,
    48'h00000400ef568,
    48'h000007b034684,
    48'h00000400ef570,
    48'h000007b034684,
    48'h00000400ef578,
    48'h000007b034684,
    48'h00000400ef580,
    48'h000007b034684,
    48'h00000400ef588,
    48'h000007b034684,
    48'h00000400ef590,
    48'h000007b034684,
    48'h00000400ef598,
    48'h000007b034684,
    48'h00000400ef5a0,
    48'h000007b034684,
    48'h00000400ef5a8,
    48'h000007b034684,
    48'h00000400ef5b0,
    48'h000007b034684,
    48'h00000400ef5b8,
    48'h000007b034684,
    48'h00000400ef5c0,
    48'h000007b034684,
    48'h00000400ef5c8,
    48'h000007b034684,
    48'h00000400ef5d0,
    48'h000007b034684,
    48'h00000400ef5d8,
    48'h000007b034684,
    48'h00000400ef5e0,
    48'h000007b034684,
    48'h00000400ef5e8,
    48'h000007b034684,
    48'h00000400ef5f0,
    48'h000007b034684,
    48'h00000400ef5f8,
    48'h000007b034684,
    48'h00000400ef600,
    48'h000007b034684,
    48'h00000400ef608,
    48'h000007b034684,
    48'h00000400ef610,
    48'h000007b034684,
    48'h00000400ef618,
    48'h000007b034684,
    48'h00000400ef620,
    48'h000007b034684,
    48'h00000400ef628,
    48'h000007b034684,
    48'h00000400ef630,
    48'h000007b034684,
    48'h00000400ef638,
    48'h000007b034684,
    48'h00000400ef640,
    48'h000007b034684,
    48'h00000400ef648,
    48'h000007b034684,
    48'h00000400ef650,
    48'h000007b034684,
    48'h00000400ef658,
    48'h000007b034684,
    48'h00000400ef660,
    48'h000007b034684,
    48'h00000400ef668,
    48'h000007b034684,
    48'h00000400ef670,
    48'h000007b034684,
    48'h00000400ef678,
    48'h000007b034684,
    48'h00000400ef680,
    48'h000007b034684,
    48'h00000400ef688,
    48'h000007b034684,
    48'h00000400ef690,
    48'h000007b034684,
    48'h00000400ef698,
    48'h000007b034684,
    48'h00000400ef6a0,
    48'h000007b034684,
    48'h00000400ef6a8,
    48'h000007b034684,
    48'h00000400ef6b0,
    48'h000007b034684,
    48'h00000400ef6b8,
    48'h000007b034684,
    48'h00000400ef6c0,
    48'h000007b034684,
    48'h00000400ef6c8,
    48'h000007b034684,
    48'h00000400ef6d0,
    48'h000007b034684,
    48'h00000400ef6d8,
    48'h000007b034684,
    48'h00000400ef6e0,
    48'h000007b034684,
    48'h00000400ef6e8,
    48'h000007b034684,
    48'h00000400ef6f0,
    48'h000007b034684,
    48'h00000400ef6f8,
    48'h000007b034684,
    48'h00000400ef700,
    48'h000007b034684,
    48'h00000400ef708,
    48'h000007b034684,
    48'h00000400ef710,
    48'h000007b034684,
    48'h00000400ef718,
    48'h000007b034684,
    48'h00000400ef720,
    48'h000007b034684,
    48'h00000400ef728,
    48'h000007b034684,
    48'h00000400ef730,
    48'h000007b034684,
    48'h00000400ef738,
    48'h000007b034684,
    48'h00000400ef740,
    48'h000007b034684,
    48'h00000400ef748,
    48'h000007b034684,
    48'h00000400ef750,
    48'h000007b034684,
    48'h00000400ef758,
    48'h000007b034684,
    48'h00000400ef760,
    48'h000007b034684,
    48'h00000400ef768,
    48'h000007b034684,
    48'h00000400ef770,
    48'h000007b034684,
    48'h00000400ef778,
    48'h000007b034684,
    48'h00000400ef780,
    48'h000007b034684,
    48'h00000400ef788,
    48'h000007b034684,
    48'h00000400ef790,
    48'h000007b034684,
    48'h00000400ef798,
    48'h000007b034684,
    48'h00000400ef7a0,
    48'h000007b034684,
    48'h00000400ef7a8,
    48'h000007b034684,
    48'h00000400ef7b0,
    48'h000007b034684,
    48'h00000400ef7b8,
    48'h000007b034684,
    48'h00000400ef7c0,
    48'h000007b034684,
    48'h00000400ef7c8,
    48'h000007b034684,
    48'h00000400ef7d0,
    48'h000007b034684,
    48'h00000400ef7d8,
    48'h000007b034684,
    48'h00000400ef7e0,
    48'h000007b034684,
    48'h00000400ef7e8,
    48'h000007b034684,
    48'h00000400ef7f0,
    48'h000007b034684,
    48'h00000400ef7f8,
    48'h000007b034684,
    48'h00000400ef800,
    48'h000007b034684,
    48'h00000400ef808,
    48'h000007b034684,
    48'h00000400ef810,
    48'h000007b034684,
    48'h00000400ef818,
    48'h000007b034684,
    48'h00000400ef820,
    48'h000007b034684,
    48'h00000400ef828,
    48'h000007b034684,
    48'h00000400ef830,
    48'h000007b034684,
    48'h00000400ef838,
    48'h000007b034684,
    48'h00000400ef840,
    48'h000007b034684,
    48'h00000400ef848,
    48'h000007b034684,
    48'h00000400ef850,
    48'h000007b034684,
    48'h00000400ef858,
    48'h000007b034684,
    48'h00000400ef860,
    48'h000007b034684,
    48'h00000400ef868,
    48'h000007b034684,
    48'h00000400ef870,
    48'h000007b034684,
    48'h00000400ef878,
    48'h000007b034684,
    48'h00000400ef880,
    48'h000007b034684,
    48'h00000400ef888,
    48'h000007b034684,
    48'h00000400ef890,
    48'h000007b034684,
    48'h00000400ef898,
    48'h000007b034684,
    48'h00000400ef8a0,
    48'h000007b034684,
    48'h00000400ef8a8,
    48'h000007b034684,
    48'h00000400ef8b0,
    48'h000007b034684,
    48'h00000400ef8b8,
    48'h000007b034684,
    48'h00000400ef8c0,
    48'h000007b034684,
    48'h00000400ef8c8,
    48'h000007b034684,
    48'h00000400ef8d0,
    48'h000007b034684,
    48'h00000400ef8d8,
    48'h000007b034684,
    48'h00000400ef8e0,
    48'h000007b034684,
    48'h00000400ef8e8,
    48'h000007b034684,
    48'h00000400ef8f0,
    48'h000007b034684,
    48'h00000400ef8f8,
    48'h000007b034684,
    48'h00000400ef900,
    48'h000007b034684,
    48'h00000400ef908,
    48'h000007b034684,
    48'h00000400ef910,
    48'h000007b034684,
    48'h00000400ef918,
    48'h000007b034684,
    48'h00000400ef920,
    48'h000007b034684,
    48'h00000400ef928,
    48'h000007b034684,
    48'h00000400ef930,
    48'h000007b034684,
    48'h00000400ef938,
    48'h000007b034684,
    48'h00000400ef940,
    48'h000007b034684,
    48'h00000400ef948,
    48'h000007b034684,
    48'h00000400ef950,
    48'h000007b034684,
    48'h00000400ef958,
    48'h000007b034684,
    48'h00000400ef960,
    48'h000007b034684,
    48'h00000400ef968,
    48'h000007b034684,
    48'h00000400ef970,
    48'h000007b034684,
    48'h00000400ef978,
    48'h000007b034684,
    48'h00000400ef980,
    48'h000007b034684,
    48'h00000400ef988,
    48'h000007b034684,
    48'h00000400ef990,
    48'h000007b034684,
    48'h00000400ef998,
    48'h000007b034684,
    48'h00000400ef9a0,
    48'h000007b034684,
    48'h00000400ef9a8,
    48'h000007b034684,
    48'h00000400ef9b0,
    48'h000007b034684,
    48'h00000400ef9b8,
    48'h000007b034684,
    48'h00000400ef9c0,
    48'h000007b034684,
    48'h00000400ef9c8,
    48'h000007b034684,
    48'h00000400ef9d0,
    48'h000007b034684,
    48'h00000400ef9d8,
    48'h000007b034684,
    48'h00000400ef9e0,
    48'h000007b034684,
    48'h00000400ef9e8,
    48'h000007b034684,
    48'h00000400ef9f0,
    48'h000007b034684,
    48'h00000400ef9f8,
    48'h000007b034684,
    48'h00000400efa00,
    48'h000007b034684,
    48'h00000400efa08,
    48'h000007b034684,
    48'h00000400efa10,
    48'h000007b034684,
    48'h00000400efa18,
    48'h000007b034684,
    48'h00000400efa20,
    48'h000007b034684,
    48'h00000400efa28,
    48'h000007b034684,
    48'h00000400efa30,
    48'h000007b034684,
    48'h00000400efa38,
    48'h000007b034684,
    48'h00000400efa40,
    48'h000007b034684,
    48'h00000400efa48,
    48'h000007b034684,
    48'h00000400efa50,
    48'h000007b034684,
    48'h00000400efa58,
    48'h000007b034684,
    48'h00000400efa60,
    48'h000007b034684,
    48'h00000400efa68,
    48'h000007b034684,
    48'h00000400efa70,
    48'h000007b034684,
    48'h00000400efa78,
    48'h000007b034684,
    48'h00000400efa80,
    48'h000007b034684,
    48'h00000400efa88,
    48'h000007b034684,
    48'h00000400efa90,
    48'h000007b034684,
    48'h00000400efa98,
    48'h000007b034684,
    48'h00000400efaa0,
    48'h000007b034684,
    48'h00000400efaa8,
    48'h000007b034684,
    48'h00000400efab0,
    48'h000007b034684,
    48'h00000400efab8,
    48'h000007b034684,
    48'h00000400efac0,
    48'h000007b034684,
    48'h00000400efac8,
    48'h000007b034684,
    48'h00000400efad0,
    48'h000007b034684,
    48'h00000400efad8,
    48'h000007b034684,
    48'h00000400efae0,
    48'h000007b034684,
    48'h00000400efae8,
    48'h000007b034684,
    48'h00000400efaf0,
    48'h000007b034684,
    48'h00000400efaf8,
    48'h000007b034684,
    48'h00000400efb00,
    48'h000007b034684,
    48'h00000400efb08,
    48'h000007b034684,
    48'h00000400efb10,
    48'h000007b034684,
    48'h00000400efb18,
    48'h000007b034684,
    48'h00000400efb20,
    48'h000007b034684,
    48'h00000400efb28,
    48'h000007b034684,
    48'h00000400efb30,
    48'h000007b034684,
    48'h00000400efb38,
    48'h000007b034684,
    48'h00000400efb40,
    48'h000007b034684,
    48'h00000400efb48,
    48'h000007b034684,
    48'h00000400efb50,
    48'h000007b034684,
    48'h00000400efb58,
    48'h000007b034684,
    48'h00000400efb60,
    48'h000007b034684,
    48'h00000400efb68,
    48'h000007b034684,
    48'h00000400efb70,
    48'h000007b034684,
    48'h00000400efb78,
    48'h000007b034684,
    48'h00000400efb80,
    48'h000007b034684,
    48'h00000400efb88,
    48'h000007b034684,
    48'h00000400efb90,
    48'h000007b034684,
    48'h00000400efb98,
    48'h000007b034684,
    48'h00000400efba0,
    48'h000007b034684,
    48'h00000400efba8,
    48'h000007b034684,
    48'h00000400efbb0,
    48'h000007b034684,
    48'h00000400efbb8,
    48'h000007b034684,
    48'h00000400efbc0,
    48'h000007b034684,
    48'h00000400efbc8,
    48'h000007b034684,
    48'h00000400efbd0,
    48'h000007b034684,
    48'h00000400efbd8,
    48'h000007b034684,
    48'h00000400efbe0,
    48'h000007b034684,
    48'h00000400efbe8,
    48'h000007b034684,
    48'h00000400efbf0,
    48'h000007b034684,
    48'h00000400efbf8,
    48'h000007b034684,
    48'h00000400efc00,
    48'h000007b034684,
    48'h00000400efc08,
    48'h000007b034684,
    48'h00000400efc10,
    48'h000007b034684,
    48'h00000400efc18,
    48'h000007b034684,
    48'h00000400efc20,
    48'h000007b034684,
    48'h00000400efc28,
    48'h000007b034684,
    48'h00000400efc30,
    48'h000007b034684,
    48'h00000400efc38,
    48'h000007b034684,
    48'h00000400efc40,
    48'h000007b034684,
    48'h00000400efc48,
    48'h000007b034684,
    48'h00000400efc50,
    48'h000007b034684,
    48'h00000400efc58,
    48'h000007b034684,
    48'h00000400efc60,
    48'h000007b034684,
    48'h00000400efc68,
    48'h000007b034684,
    48'h00000400efc70,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b0337fc,
    48'h00000400e5414,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c08,
    48'h00000400321e8,
    48'h0000040032338,
    48'h00000400ed254,
    48'h00000400ed25c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03473c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032338,
    48'h00000400ed274,
    48'h00000400ed274,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034534,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003234c,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020474,
    48'h0000040020474,
    48'h00000400e53f4,
    48'h000007b0337fc,
    48'h00000400e53c8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h00000400edc98,
    48'h000007b034400,
    48'h00000400edc9c,
    48'h000007b034404,
    48'h000007b034400,
    48'h000007b034404,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034400,
    48'h000007b034404,
    48'h000007b03447c,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b034514,
    48'h000007b034510,
    48'h0000040059780,
    48'h000007b034404,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073d04,
    48'h000007b034510,
    48'h0000040073d04,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034510,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040097014,
    48'h000007b034538,
    48'h0000040097014,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h000007b034538,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0345cc,
    48'h000007b0345cc,
    48'h0000040020544,
    48'h000007b03464c,
    48'h000007b03464c,
    48'h000007b0346c4,
    48'h0000040020054,
    48'h000007b0346c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0345c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h000007b034400,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h000007b034400,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000007b034400,
    48'h000004003bfb8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345c4,
    48'h000007b034514,
    48'h000007b0345c4,
    48'h000007b0345c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000007b034400,
    48'h0000040032350,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034538,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b034514,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h000007b034404,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073d04,
    48'h000007b0345fc,
    48'h0000040073d04,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0345fc,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034514,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034514,
    48'h00000400efc84,
    48'h00000400efc88,
    48'h000007b034400,
    48'h0000040020468,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfb8,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfb8,
    48'h00000400efc90,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c20,
    48'h0000040045c20,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020614,
    48'h0000040020344,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b0344fc,
    48'h0000040020610,
    48'h0000040020614,
    48'h000004000e43c,
    48'h000007b0344fc,
    48'h000007b0344fc,
    48'h0000040059918,
    48'h000007b0337fc,
    48'h000007b0344fc,
    48'h00000400597c0,
    48'h0000040020610,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b034504,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b034504,
    48'h000007b0345b0,
    48'h000007b0345ac,
    48'h000007b0345a8,
    48'h0000040020614,
    48'h000004000e43c,
    48'h000007b0345b4,
    48'h000007b0345b4,
    48'h0000040059914,
    48'h00000400d602c,
    48'h000007b0345b0,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e5434,
    48'h00000400e53e8,
    48'h00000400e53e4,
    48'h000007b0345b4,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345c4,
    48'h000007b0345c0,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345c4,
    48'h000007b0345c0,
    48'h000007b03467c,
    48'h000007b034678,
    48'h000007b034674,
    48'h000007b034670,
    48'h0000040020748,
    48'h000007b03466c,
    48'h0000040058f58,
    48'h000007b03466c,
    48'h000007b034668,
    48'h000007b0345a8,
    48'h00000400e5400,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b03470c,
    48'h000007b034708,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf4,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6aac,
    48'h00000400e6ab4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6acc,
    48'h000007b0345ac,
    48'h00000400e6acc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345ac,
    48'h000007b03468c,
    48'h000007b03468c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003234c,
    48'h000007b0345a8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345a8,
    48'h00000400e53fc,
    48'h000007b0337fc,
    48'h0000040020470,
    48'h0000040020470,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e53e4,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e5408,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b03463c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70c0,
    48'h000007b03464c,
    48'h000007b034648,
    48'h000007b034644,
    48'h000007b03464c,
    48'h000007b034648,
    48'h000007b034644,
    48'h000007b0337fc,
    48'h000007b03463c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bfc,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70bc,
    48'h00000400e70c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70d8,
    48'h00000400e70d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345b0,
    48'h00000400e53e0,
    48'h000007b0345a8,
    48'h000007b034400,
    48'h00000400edc98,
    48'h000007b034404,
    48'h00000400edc9c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004002078c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032350,
    48'h000004002062c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h000004002079c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03438c,
    48'h000007b03438c,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h000007b03447c,
    48'h000004002078c,
    48'h0000040020618,
    48'h000007b0337fc,
    48'h000004002061c,
    48'h000004000e43c,
    48'h000007b03447c,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b034534,
    48'h0000040020618,
    48'h000004002061c,
    48'h000004000e43c,
    48'h000007b03453c,
    48'h000007b03453c,
    48'h0000040059918,
    48'h000007b0337fc,
    48'h0000040020618,
    48'h00000400e5434,
    48'h00000400e53e8,
    48'h000007b03453c,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b0345f8,
    48'h000007b0345f4,
    48'h000007b0345f0,
    48'h0000040020748,
    48'h000007b0345ec,
    48'h0000040058f58,
    48'h000007b0345ec,
    48'h000007b0345e8,
    48'h000007b034538,
    48'h00000400e5400,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf4,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6aac,
    48'h00000400e6ab4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6acc,
    48'h000007b034534,
    48'h00000400e6acc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034534,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003234c,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h00000400e53fc,
    48'h000007b0337fc,
    48'h0000040020470,
    48'h0000040020470,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h00000400edca0,
    48'h000007b034400,
    48'h00000400edca4,
    48'h000007b034404,
    48'h000007b034400,
    48'h000007b034404,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034400,
    48'h000007b034404,
    48'h000007b03447c,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b034514,
    48'h000007b034510,
    48'h0000040059780,
    48'h000007b034404,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073d08,
    48'h000007b034510,
    48'h0000040073d08,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034510,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040097018,
    48'h000007b034538,
    48'h0000040097018,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h000007b034538,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0345cc,
    48'h000007b0345cc,
    48'h0000040020544,
    48'h000007b03464c,
    48'h000007b03464c,
    48'h000007b0346c4,
    48'h0000040020054,
    48'h000007b0346c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0345c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h000007b034400,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h000007b034400,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000007b034400,
    48'h000004003bfbc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345c4,
    48'h000007b034514,
    48'h000007b0345c4,
    48'h000007b0345c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000007b034400,
    48'h0000040032354,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034538,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b034514,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h000007b034404,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073d08,
    48'h000007b0345fc,
    48'h0000040073d08,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0345fc,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034514,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034514,
    48'h00000400f014c,
    48'h00000400f0150,
    48'h000007b034400,
    48'h0000040020468,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfbc,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfbc,
    48'h00000400f0158,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c24,
    48'h0000040045c24,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004002061c,
    48'h0000040020344,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b0344fc,
    48'h0000040020618,
    48'h000004002061c,
    48'h000004000e43c,
    48'h000007b0344fc,
    48'h000007b0344fc,
    48'h0000040059918,
    48'h000007b0337fc,
    48'h000007b0344fc,
    48'h00000400597c0,
    48'h0000040020618,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b034504,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b034504,
    48'h000007b0345b0,
    48'h000007b0345ac,
    48'h000007b0345a8,
    48'h000004002061c,
    48'h000004000e43c,
    48'h000007b0345b4,
    48'h000007b0345b4,
    48'h0000040059914,
    48'h00000400d602c,
    48'h000007b0345b0,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e5434,
    48'h00000400e53e8,
    48'h00000400e53e4,
    48'h000007b0345b4,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345c4,
    48'h000007b0345c0,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345c4,
    48'h000007b0345c0,
    48'h000007b03467c,
    48'h000007b034678,
    48'h000007b034674,
    48'h000007b034670,
    48'h0000040020748,
    48'h000007b03466c,
    48'h0000040058f58,
    48'h000007b03466c,
    48'h000007b034668,
    48'h000007b0345a8,
    48'h00000400e5400,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b03470c,
    48'h000007b034708,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf4,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6aac,
    48'h00000400e6ab4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6acc,
    48'h000007b0345ac,
    48'h00000400e6acc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345ac,
    48'h000007b03468c,
    48'h000007b03468c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003234c,
    48'h000007b0345a8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345a8,
    48'h00000400e53fc,
    48'h000007b0337fc,
    48'h0000040020470,
    48'h0000040020470,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e53e4,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e5408,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b03463c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70c0,
    48'h000007b03464c,
    48'h000007b034648,
    48'h000007b034644,
    48'h000007b03464c,
    48'h000007b034648,
    48'h000007b034644,
    48'h000007b0337fc,
    48'h000007b03463c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bfc,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70bc,
    48'h00000400e70c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70d8,
    48'h00000400e70d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345b0,
    48'h00000400e53e0,
    48'h000007b0345a8,
    48'h000007b034400,
    48'h00000400edca0,
    48'h000007b034404,
    48'h00000400edca4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004002078c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032354,
    48'h0000040020630,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h000004002079c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03438c,
    48'h000007b03438c,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h000007b03447c,
    48'h000004002078c,
    48'h0000040020620,
    48'h000007b0337fc,
    48'h0000040020624,
    48'h000004000e43c,
    48'h000007b03447c,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b034534,
    48'h0000040020620,
    48'h0000040020624,
    48'h000004000e43c,
    48'h000007b03453c,
    48'h000007b03453c,
    48'h0000040059918,
    48'h000007b0337fc,
    48'h0000040020620,
    48'h00000400e5434,
    48'h00000400e53e8,
    48'h000007b03453c,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b0345f8,
    48'h000007b0345f4,
    48'h000007b0345f0,
    48'h0000040020748,
    48'h000007b0345ec,
    48'h0000040058f58,
    48'h000007b0345ec,
    48'h000007b0345e8,
    48'h000007b034538,
    48'h00000400e5400,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf4,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6aac,
    48'h00000400e6ab4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6acc,
    48'h000007b034534,
    48'h00000400e6acc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034534,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003234c,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h00000400e53fc,
    48'h000007b0337fc,
    48'h0000040020470,
    48'h0000040020470,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h00000400edca8,
    48'h000007b034400,
    48'h00000400edcac,
    48'h000007b034404,
    48'h000007b034400,
    48'h000007b034404,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034400,
    48'h000007b034404,
    48'h000007b03447c,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b034514,
    48'h000007b034510,
    48'h0000040059780,
    48'h000007b034404,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073d0c,
    48'h000007b034510,
    48'h0000040073d0c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034510,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h000004009701c,
    48'h000007b034538,
    48'h000004009701c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h000007b034538,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0345cc,
    48'h000007b0345cc,
    48'h0000040020544,
    48'h000007b03464c,
    48'h000007b03464c,
    48'h000007b0346c4,
    48'h0000040020054,
    48'h000007b0346c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0345c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h000007b034400,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h000007b034400,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000007b034400,
    48'h000004003bfc0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345c4,
    48'h000007b034514,
    48'h000007b0345c4,
    48'h000007b0345c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000007b034400,
    48'h0000040032358,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034538,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b034514,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h000007b034404,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073d0c,
    48'h000007b0345fc,
    48'h0000040073d0c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0345fc,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034514,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034514,
    48'h00000400f0614,
    48'h00000400f0618,
    48'h000007b034400,
    48'h0000040020468,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfc0,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfc0,
    48'h00000400f0620,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c28,
    48'h0000040045c28,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020624,
    48'h0000040020344,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b0344fc,
    48'h0000040020620,
    48'h0000040020624,
    48'h000004000e43c,
    48'h000007b0344fc,
    48'h000007b0344fc,
    48'h0000040059918,
    48'h000007b0337fc,
    48'h000007b0344fc,
    48'h00000400597c0,
    48'h0000040020620,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b034504,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b034504,
    48'h000007b0345b0,
    48'h000007b0345ac,
    48'h000007b0345a8,
    48'h0000040020624,
    48'h000004000e43c,
    48'h000007b0345b4,
    48'h000007b0345b4,
    48'h0000040059914,
    48'h00000400d602c,
    48'h000007b0345b0,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e5434,
    48'h00000400e53e8,
    48'h00000400e53e4,
    48'h000007b0345b4,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345c4,
    48'h000007b0345c0,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345c4,
    48'h000007b0345c0,
    48'h000007b03467c,
    48'h000007b034678,
    48'h000007b034674,
    48'h000007b034670,
    48'h0000040020748,
    48'h000007b03466c,
    48'h0000040058f58,
    48'h000007b03466c,
    48'h000007b034668,
    48'h000007b0345a8,
    48'h00000400e5400,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b03470c,
    48'h000007b034708,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bf4,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6aac,
    48'h00000400e6ab4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032324,
    48'h00000400e6acc,
    48'h000007b0345ac,
    48'h00000400e6acc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345ac,
    48'h000007b03468c,
    48'h000007b03468c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003234c,
    48'h000007b0345a8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345a8,
    48'h00000400e53fc,
    48'h000007b0337fc,
    48'h0000040020470,
    48'h0000040020470,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e53e4,
    48'h000007b0337fc,
    48'h000007b0345b0,
    48'h00000400e5408,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b03463c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70c0,
    48'h000007b03464c,
    48'h000007b034648,
    48'h000007b034644,
    48'h000007b03464c,
    48'h000007b034648,
    48'h000007b034644,
    48'h000007b0337fc,
    48'h000007b03463c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045bfc,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70bc,
    48'h00000400e70c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003232c,
    48'h00000400e70d8,
    48'h00000400e70d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345b0,
    48'h00000400e53e0,
    48'h000007b0345a8,
    48'h000007b034400,
    48'h00000400edca8,
    48'h000007b034404,
    48'h00000400edcac,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004002078c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032358,
    48'h0000040020634,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h000004002079c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004002035c,
    48'h000004002034c,
    48'h0000040020354,
    48'h0000040020350,
    48'h0000040020358,
    48'h0000040020350,
    48'h000004002035a,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004002035c,
    48'h000007b03438c,
    48'h000007b03438c,
    48'h000007b034404,
    48'h000007b034400,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b0344e8,
    48'h0000040020358,
    48'h000004002048e,
    48'h000004000e43c,
    48'h000007b034484,
    48'h0000040020358,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034484,
    48'h0000040020354,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b03448c,
    48'h000007b034488,
    48'h0000040020438,
    48'h000007b0337fc,
    48'h00000400597d0,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b03458c,
    48'h000007b034588,
    48'h000007b03458c,
    48'h000007b034588,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b40,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b974,
    48'h000004005b97c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b994,
    48'h0000040020438,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020438,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020358,
    48'h000004000e43c,
    48'h000007b034400,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b0344bc,
    48'h000007b0344b8,
    48'h000007b0344b4,
    48'h000007b0344b0,
    48'h0000040020354,
    48'h0000040020358,
    48'h000004000e43c,
    48'h000007b0344bc,
    48'h000007b0344bc,
    48'h00000400597f8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b58,
    48'h00000400321e8,
    48'h0000040032288,
    48'h00000400ba2e4,
    48'h00000400ba2ec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032288,
    48'h00000400ba304,
    48'h000007b0344b8,
    48'h00000400ba304,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0344b8,
    48'h000007b0337fc,
    48'h000007b0344b8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b034540,
    48'h0000040020358,
    48'h000004000e43c,
    48'h000007b034544,
    48'h000007b034544,
    48'h0000040059830,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b90,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6154,
    48'h00000400d615c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6170,
    48'h000007b0344b4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0344b4,
    48'h000007b034544,
    48'h000004005983c,
    48'h0000040059838,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b88,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b44,
    48'h00000400d5b4c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b60,
    48'h000007b034540,
    48'h00000400d5b60,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h00000400207cc,
    48'h000004002077c,
    48'h00000400207bc,
    48'h000007b0345fc,
    48'h000007b0345f8,
    48'h000007b0345f4,
    48'h000007b0345f0,
    48'h0000040020790,
    48'h00000400207cc,
    48'h0000040020358,
    48'h0000040020068,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h000007b034668,
    48'h0000040020358,
    48'h000004002048e,
    48'h000004000e43c,
    48'h000007b0345f4,
    48'h0000040020358,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f4,
    48'h0000040059838,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b4c,
    48'h000007b0345fc,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345fc,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h0000040059838,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b88,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b44,
    48'h00000400d5b4c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b60,
    48'h000007b0345f8,
    48'h00000400d5b60,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f8,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h0000040059770,
    48'h000007b0337fc,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h000007b034684,
    48'h0000040020054,
    48'h000007b034684,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0344b4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f4,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b0346bc,
    48'h000007b0344b4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h000007b0345f8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761d4,
    48'h000007b0346bc,
    48'h00000400761d4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0346bc,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0346b4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0344b4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b0344b4,
    48'h00000400f0bc8,
    48'h000007b0344b4,
    48'h00000400f0be0,
    48'h000007b0344b4,
    48'h00000400f0be8,
    48'h000007b0344b4,
    48'h00000400f0bf4,
    48'h000007b0344b4,
    48'h00000400f0bfc,
    48'h000007b0344b4,
    48'h00000400f0c08,
    48'h000007b0344b4,
    48'h00000400f0c14,
    48'h000007b0344b4,
    48'h00000400f0c20,
    48'h000007b0344b4,
    48'h00000400f0b08,
    48'h0000040020730,
    48'h000007b0344b4,
    48'h00000400f0b0c,
    48'h000007b0344b4,
    48'h00000400f0ae0,
    48'h000007b0344b4,
    48'h00000400f0bd4,
    48'h000007b0344b4,
    48'h00000400f0b10,
    48'h000007b0344b4,
    48'h00000400f0b28,
    48'h000007b0344b4,
    48'h00000400f0b14,
    48'h000007b0344b4,
    48'h00000400f0b1c,
    48'h000007b0344b4,
    48'h00000400f0c2c,
    48'h000007b0344b4,
    48'h00000400f0b34,
    48'h000007b0344b4,
    48'h00000400f0b6c,
    48'h000007b0337fc,
    48'h000007b0344b4,
    48'h0000040020068,
    48'h000007b0345f4,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03467c,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0347fc,
    48'h000007b0347f8,
    48'h000007b0347d4,
    48'h000007b0347d0,
    48'h0000040059780,
    48'h00000400f0b38,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761c4,
    48'h000007b0347d0,
    48'h00000400761c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b0347d0,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994d4,
    48'h000007b0347f8,
    48'h00000400994d4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b34,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034884,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h0000040020544,
    48'h000007b03490c,
    48'h000007b03490c,
    48'h000007b034984,
    48'h0000040020054,
    48'h000007b034984,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034884,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b34,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b34,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b34,
    48'h000004003bfc4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034884,
    48'h000007b0347d4,
    48'h000007b034884,
    48'h000007b034884,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b34,
    48'h000004003235c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b0348bc,
    48'h000007b0347d4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0b38,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761c4,
    48'h000007b0348bc,
    48'h00000400761c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0348bc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0348b4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0347d4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347d4,
    48'h00000400f0c64,
    48'h00000400f0c68,
    48'h00000400f0b34,
    48'h0000040020468,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfc4,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfc4,
    48'h00000400f0c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c2c,
    48'h0000040045c2c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347f8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0347fc,
    48'h000007b0347f8,
    48'h000007b0347d4,
    48'h000007b0347d0,
    48'h0000040059780,
    48'h00000400f0b2c,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761d0,
    48'h000007b0347d0,
    48'h00000400761d0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b0347d0,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994e0,
    48'h000007b0347f8,
    48'h00000400994e0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b28,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034884,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h0000040020544,
    48'h000007b03490c,
    48'h000007b03490c,
    48'h000007b034984,
    48'h0000040020054,
    48'h000007b034984,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034884,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b28,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b28,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b28,
    48'h000004003bfc8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034884,
    48'h000007b0347d4,
    48'h000007b034884,
    48'h000007b034884,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b28,
    48'h0000040032360,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b0348bc,
    48'h000007b0347d4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0b2c,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761d0,
    48'h000007b0348bc,
    48'h00000400761d0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0348bc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0348b4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0347d4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347d4,
    48'h00000400f0cac,
    48'h00000400f0cb0,
    48'h00000400f0b28,
    48'h0000040020468,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfc8,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfc8,
    48'h00000400f0cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h0000040045c30,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347f8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h00000400f0b70,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0347fc,
    48'h000007b0347f8,
    48'h000007b0347d4,
    48'h000007b0347d0,
    48'h0000040059780,
    48'h00000400f0b70,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761cc,
    48'h000007b0347d0,
    48'h00000400761cc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b0347d0,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994dc,
    48'h000007b0347f8,
    48'h00000400994dc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b6c,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034884,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h0000040020544,
    48'h000007b03490c,
    48'h000007b03490c,
    48'h000007b034984,
    48'h0000040020054,
    48'h000007b034984,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034884,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b6c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b6c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b6c,
    48'h000004003bfcc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034884,
    48'h000007b0347d4,
    48'h000007b034884,
    48'h000007b034884,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b6c,
    48'h0000040032364,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b0348bc,
    48'h000007b0347d4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0b70,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761cc,
    48'h000007b0348bc,
    48'h00000400761cc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0348bc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0348b4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0347d4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347d4,
    48'h00000400f0cf4,
    48'h00000400f0cf8,
    48'h00000400f0b6c,
    48'h0000040020468,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfcc,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfcc,
    48'h00000400f0d00,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c34,
    48'h0000040045c34,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347f8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b6c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032364,
    48'h00000400f0b9c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400f0b7c,
    48'h000007b0337fc,
    48'h00000400f0b28,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cac,
    48'h000007b034724,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cb0,
    48'h000007b034728,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cb4,
    48'h000007b03472c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cb8,
    48'h000007b034730,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cbc,
    48'h000007b034734,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cc0,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h00000400f0af8,
    48'h00000400f0b44,
    48'h000007b0337fc,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b10,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b10,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b10,
    48'h000004003bfd0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b10,
    48'h0000040032368,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b10,
    48'h0000040032368,
    48'h00000400f0d40,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b10,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d3c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d50,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d4c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d44,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfd0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c38,
    48'h0000040045c38,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c38,
    48'h0000040045c38,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c38,
    48'h0000040045c38,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c38,
    48'h0000040045c38,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c38,
    48'h0000040045c38,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c38,
    48'h0000040045c38,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d38,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d3c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b10,
    48'h0000040045c38,
    48'h0000040045c38,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b10,
    48'h0000040045c38,
    48'h0000040045c38,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b10,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d44,
    48'h00000400f0d44,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d40,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b14,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b14,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b14,
    48'h000004003bfd4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b14,
    48'h000004003236c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b14,
    48'h000004003236c,
    48'h00000400f0d88,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b14,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d84,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d98,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d94,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d8c,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfd4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c3c,
    48'h0000040045c3c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c3c,
    48'h0000040045c3c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c3c,
    48'h0000040045c3c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c3c,
    48'h0000040045c3c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c3c,
    48'h0000040045c3c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c3c,
    48'h0000040045c3c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d80,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d84,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b14,
    48'h0000040045c3c,
    48'h0000040045c3c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b14,
    48'h0000040045c3c,
    48'h0000040045c3c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b14,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d8c,
    48'h00000400f0d8c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d88,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347bc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b034838,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b034838,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b034944,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h0000040020544,
    48'h000007b0349cc,
    48'h000007b0349cc,
    48'h000007b034a44,
    48'h0000040020054,
    48'h000007b034a44,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034944,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b18,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b18,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b18,
    48'h000004003bfd8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034944,
    48'h000007b034944,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b18,
    48'h0000040032370,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b18,
    48'h0000040032370,
    48'h00000400f0dd0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b18,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348c0,
    48'h000007b0348bc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348c0,
    48'h000007b0348bc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0dcc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0de0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0ddc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0dd4,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfd8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c40,
    48'h0000040045c40,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c40,
    48'h0000040045c40,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c40,
    48'h0000040045c40,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c40,
    48'h0000040045c40,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c40,
    48'h0000040045c40,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c40,
    48'h0000040045c40,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0dc8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0dcc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b18,
    48'h0000040045c40,
    48'h0000040045c40,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b18,
    48'h0000040045c40,
    48'h0000040045c40,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b18,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0dd4,
    48'h00000400f0dd4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0dd0,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b18,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h000007b0347bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b1c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b1c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b1c,
    48'h000004003bfdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b1c,
    48'h0000040032374,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b1c,
    48'h0000040032374,
    48'h00000400f0e18,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b1c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0e14,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0e28,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0e24,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0e1c,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfdc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c44,
    48'h0000040045c44,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c44,
    48'h0000040045c44,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c44,
    48'h0000040045c44,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c44,
    48'h0000040045c44,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c44,
    48'h0000040045c44,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c44,
    48'h0000040045c44,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0e10,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0e14,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b1c,
    48'h0000040045c44,
    48'h0000040045c44,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b1c,
    48'h0000040045c44,
    48'h0000040045c44,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b1c,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0e1c,
    48'h00000400f0e1c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0e18,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b1c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032374,
    48'h00000400f0b88,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b20,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b20,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b20,
    48'h000004003bfe0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b20,
    48'h0000040032378,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b20,
    48'h0000040032378,
    48'h00000400f0e60,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b20,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0e5c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0e70,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0e6c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0e64,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfe0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c48,
    48'h0000040045c48,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c48,
    48'h0000040045c48,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c48,
    48'h0000040045c48,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c48,
    48'h0000040045c48,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c48,
    48'h0000040045c48,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c48,
    48'h0000040045c48,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0e58,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0e5c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b20,
    48'h0000040045c48,
    48'h0000040045c48,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b20,
    48'h0000040045c48,
    48'h0000040045c48,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b20,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0e64,
    48'h00000400f0e64,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0e60,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b20,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032378,
    48'h00000400f0b8c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b24,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b24,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b24,
    48'h000004003bfe4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b24,
    48'h000004003237c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b24,
    48'h000004003237c,
    48'h00000400f0ea8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b24,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0ea4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0eb8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0eb4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0eac,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfe4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c4c,
    48'h0000040045c4c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c4c,
    48'h0000040045c4c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c4c,
    48'h0000040045c4c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c4c,
    48'h0000040045c4c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c4c,
    48'h0000040045c4c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c4c,
    48'h0000040045c4c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0ea0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0ea4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b24,
    48'h0000040045c4c,
    48'h0000040045c4c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b24,
    48'h0000040045c4c,
    48'h0000040045c4c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b24,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0eac,
    48'h00000400f0eac,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0ea8,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b24,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003237c,
    48'h00000400f0b90,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b54,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b5c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b5c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b5c,
    48'h000004003bfe8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b5c,
    48'h0000040032380,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b5c,
    48'h0000040032380,
    48'h00000400f0ef0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b5c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0eec,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0f00,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0efc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0ef4,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfe8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c50,
    48'h0000040045c50,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c50,
    48'h0000040045c50,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c50,
    48'h0000040045c50,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c50,
    48'h0000040045c50,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c50,
    48'h0000040045c50,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c50,
    48'h0000040045c50,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0ee8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0eec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b5c,
    48'h0000040045c50,
    48'h0000040045c50,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b5c,
    48'h0000040045c50,
    48'h0000040045c50,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b5c,
    48'h00000400f0b54,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0ef4,
    48'h00000400f0ef4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0ef0,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b5c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032380,
    48'h00000400f0b94,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b54,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0b60,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0b60,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0b60,
    48'h000004003bfec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b60,
    48'h0000040032384,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0b60,
    48'h0000040032384,
    48'h00000400f0f38,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b60,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0f34,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0f48,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0f44,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0f3c,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bfec,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c54,
    48'h0000040045c54,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c54,
    48'h0000040045c54,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c54,
    48'h0000040045c54,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c54,
    48'h0000040045c54,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c54,
    48'h0000040045c54,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c54,
    48'h0000040045c54,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0f30,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0f34,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b60,
    48'h0000040045c54,
    48'h0000040045c54,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f0b60,
    48'h0000040045c54,
    48'h0000040045c54,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b60,
    48'h00000400f0b54,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0f3c,
    48'h00000400f0f3c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0f38,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b60,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032384,
    48'h00000400f0b98,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b48,
    48'h00000400f0b64,
    48'h00000400f0b68,
    48'h00000400f0b58,
    48'h000007b0337fc,
    48'h00000400f0b44,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020344,
    48'h00000400f0b0c,
    48'h000007b0337fc,
    48'h00000400f0bcc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f0bcc,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761ac,
    48'h000007b034710,
    48'h00000400761ac,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994bc,
    48'h000007b034738,
    48'h00000400994bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0bc8,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0bc8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0bc8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0bc8,
    48'h000004003bff0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0bc8,
    48'h0000040032388,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0bcc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761ac,
    48'h000007b0347fc,
    48'h00000400761ac,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f0f7c,
    48'h00000400f0f80,
    48'h00000400f0bc8,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bff0,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bff0,
    48'h00000400f0f88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c58,
    48'h0000040045c58,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f0be4,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761b0,
    48'h000007b034710,
    48'h00000400761b0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994c0,
    48'h000007b034738,
    48'h00000400994c0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0be0,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0be0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0be0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0be0,
    48'h000004003bff4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0be0,
    48'h000004003238c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0be4,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761b0,
    48'h000007b0347fc,
    48'h00000400761b0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f0fc4,
    48'h00000400f0fc8,
    48'h00000400f0be0,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bff4,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bff4,
    48'h00000400f0fd0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c5c,
    48'h0000040045c5c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f0bec,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761b4,
    48'h000007b034710,
    48'h00000400761b4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994c4,
    48'h000007b034738,
    48'h00000400994c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0be8,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0be8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0be8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0be8,
    48'h000004003bff8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0be8,
    48'h0000040032390,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0bec,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761b4,
    48'h000007b0347fc,
    48'h00000400761b4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f194c,
    48'h00000400f1950,
    48'h00000400f0be8,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bff8,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bff8,
    48'h00000400f1958,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c60,
    48'h0000040045c60,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f0bf8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761b8,
    48'h000007b034710,
    48'h00000400761b8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994c8,
    48'h000007b034738,
    48'h00000400994c8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0bf4,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0bf4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0bf4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0bf4,
    48'h000004003bffc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0bf4,
    48'h0000040032394,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0bf8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761b8,
    48'h000007b0347fc,
    48'h00000400761b8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f22d4,
    48'h00000400f22d8,
    48'h00000400f0bf4,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bffc,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003bffc,
    48'h00000400f22e0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c64,
    48'h0000040045c64,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f0c00,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761bc,
    48'h000007b034710,
    48'h00000400761bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994cc,
    48'h000007b034738,
    48'h00000400994cc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0bfc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0bfc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0bfc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0bfc,
    48'h000004003c000,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0bfc,
    48'h0000040032398,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0c00,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761bc,
    48'h000007b0347fc,
    48'h00000400761bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f241c,
    48'h00000400f2420,
    48'h00000400f0bfc,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c000,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c000,
    48'h00000400f2428,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c68,
    48'h0000040045c68,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f0c0c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761c0,
    48'h000007b034710,
    48'h00000400761c0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994d0,
    48'h000007b034738,
    48'h00000400994d0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0c08,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f0c08,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f0c08,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f0c08,
    48'h000004003c004,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f0c08,
    48'h000004003239c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f0c0c,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761c0,
    48'h000007b0347fc,
    48'h00000400761c0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f2564,
    48'h00000400f2568,
    48'h00000400f0c08,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c004,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c004,
    48'h00000400f2570,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c6c,
    48'h0000040045c6c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h00000400f0c10,
    48'h000007b0337fc,
    48'h00000400f0c1c,
    48'h000007b0337fc,
    48'h00000400f0c30,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f4,
    48'h0000040059830,
    48'h000007b0344b4,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03467c,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b0337fc,
    48'h000007b03467c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b90,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6154,
    48'h00000400d615c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03467c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6170,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000004002077c,
    48'h00000400207bc,
    48'h00000400207cc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034544,
    48'h0000040058f58,
    48'h0000040020344,
    48'h000007b0344b4,
    48'h00000400f0b0c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0344bc,
    48'h00000400597e8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b54,
    48'h00000400321e8,
    48'h0000040032284,
    48'h00000400a2b9c,
    48'h00000400a2ba4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032284,
    48'h00000400a2bbc,
    48'h000007b034404,
    48'h00000400a2bbc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0344b4,
    48'h00000400f0bd4,
    48'h000007b034404,
    48'h00000400f0af8,
    48'h000007b0337fc,
    48'h000007b0344bc,
    48'h000007b0344b4,
    48'h000007b034404,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344c4,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344c4,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h00000400f0b44,
    48'h00000400f0af8,
    48'h00000400f0b44,
    48'h00000400f0af8,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b0345f8,
    48'h000007b0345f4,
    48'h000007b0345f0,
    48'h0000040020748,
    48'h000007b0345ec,
    48'h0000040058f58,
    48'h000007b0345ec,
    48'h000007b0345e8,
    48'h000007b034538,
    48'h00000400f0b10,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c38,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d3c,
    48'h00000400f0d44,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d58,
    48'h000007b03453c,
    48'h00000400f0d58,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03453c,
    48'h00000400f0b14,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c3c,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d84,
    48'h00000400f0d8c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0da0,
    48'h000007b0345f8,
    48'h00000400f0da0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f8,
    48'h000007b0337fc,
    48'h00000400f0b28,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cac,
    48'h00000400f0cb4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cc8,
    48'h000007b0345fc,
    48'h00000400f0cc8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345fc,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b034694,
    48'h000007b034690,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h0000040059770,
    48'h000007b034698,
    48'h0000040059774,
    48'h000007b03469c,
    48'h0000040059778,
    48'h000007b0346a0,
    48'h000004005977c,
    48'h000007b0346a4,
    48'h0000040059780,
    48'h000007b0346a8,
    48'h0000040059784,
    48'h000007b0346ac,
    48'h0000040059788,
    48'h000007b0346b0,
    48'h000004005978c,
    48'h000007b0346b4,
    48'h0000040059790,
    48'h000007b0346b8,
    48'h0000040059794,
    48'h000007b0346bc,
    48'h00000400f0b28,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cb4,
    48'h000007b034694,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034694,
    48'h00000400f0b28,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c30,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cac,
    48'h00000400f0cb4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032360,
    48'h00000400f0cc8,
    48'h000007b034690,
    48'h00000400f0cc8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b03477c,
    48'h000007b034778,
    48'h000007b034754,
    48'h000007b034750,
    48'h000007b0346a8,
    48'h000007b034690,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761c8,
    48'h000007b034750,
    48'h00000400761c8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346b8,
    48'h000007b034750,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994d8,
    48'h000007b034778,
    48'h00000400994d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03453c,
    48'h000007b034778,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034804,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03480c,
    48'h000007b03480c,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h000007b034904,
    48'h0000040020054,
    48'h000007b034904,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034804,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h000007b03453c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h000007b03453c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000007b03453c,
    48'h000004003c008,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034804,
    48'h000007b034754,
    48'h000007b034804,
    48'h000007b034804,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000007b03453c,
    48'h00000400323a0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034778,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03483c,
    48'h000007b034754,
    48'h000007b0337fc,
    48'h000007b0346a8,
    48'h000007b034690,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761c8,
    48'h000007b03483c,
    48'h00000400761c8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346b4,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034834,
    48'h000007b0337fc,
    48'h000007b034698,
    48'h000007b034754,
    48'h000007b034698,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034754,
    48'h00000400f28ec,
    48'h00000400f28f0,
    48'h000007b03453c,
    48'h0000040020468,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c008,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c008,
    48'h00000400f28f8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c70,
    48'h0000040045c70,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034778,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b08,
    48'h00000400f0b04,
    48'h000007b0337fc,
    48'h00000400f0b10,
    48'h000007b03453c,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c38,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d3c,
    48'h00000400f0d44,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03473c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032368,
    48'h00000400f0d58,
    48'h00000400f0d58,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b18,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0dd0,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c40,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0dcc,
    48'h00000400f0dd4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032370,
    48'h00000400f0de8,
    48'h00000400f0de8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f0b14,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c3c,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0d84,
    48'h00000400f0d8c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03473c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003236c,
    48'h00000400f0da0,
    48'h00000400f0da0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400597c0,
    48'h00000400f0ae4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03453c,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a0,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020474,
    48'h0000040020474,
    48'h00000400f0b44,
    48'h00000400f0b04,
    48'h000007b0337fc,
    48'h00000400f0ad8,
    48'h000007b03453c,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b0346c4,
    48'h000007b0346c0,
    48'h00000400207bc,
    48'h0000040020784,
    48'h000007b0346bc,
    48'h00000400205d8,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a0,
    48'h000007b0346c0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a0,
    48'h00000400f28f4,
    48'h000007b0346c4,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346c0,
    48'h000007b0346c4,
    48'h0000040020728,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h000007b0344b0,
    48'h000007b0337fc,
    48'h00000400207f8,
    48'h000007b0337fc,
    48'h0000040020788,
    48'h0000040020790,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0344b0,
    48'h000007b0344b4,
    48'h00000400f0af0,
    48'h0000040020438,
    48'h000007b0337fc,
    48'h000004002079c,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h00000400597e0,
    48'h0000040020354,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03447c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032274,
    48'h00000400730c0,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b0337fc,
    48'h000007b03447c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b44,
    48'h00000400321e8,
    48'h0000040032274,
    48'h00000400730bc,
    48'h00000400730c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032274,
    48'h00000400730d8,
    48'h00000400730d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h00000400597d0,
    48'h0000040020354,
    48'h0000040020438,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03447c,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b0337fc,
    48'h000007b03447c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b40,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b974,
    48'h000004005b97c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03447c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b994,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000004002079c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034384,
    48'h0000040020344,
    48'h000007b034380,
    48'h000007b03437c,
    48'h000007b03438c,
    48'h000007b03438c,
    48'h000007b034404,
    48'h000007b034400,
    48'h000007b03440c,
    48'h000007b03440c,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b03448c,
    48'h000007b0344e8,
    48'h000007b034380,
    48'h000004002048e,
    48'h000004000e43c,
    48'h000007b034484,
    48'h000007b034380,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034484,
    48'h000007b03437c,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034384,
    48'h000007b0337fc,
    48'h00000400597d0,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b03458c,
    48'h000007b034588,
    48'h000007b03458c,
    48'h000007b034588,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b40,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b974,
    48'h000004005b97c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b99c,
    48'h000007b034384,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034384,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b034380,
    48'h000004000e43c,
    48'h000007b034400,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b0344bc,
    48'h000007b0344b8,
    48'h000007b0344b4,
    48'h000007b0344b0,
    48'h000007b03437c,
    48'h000007b034380,
    48'h000004000e43c,
    48'h000007b0344bc,
    48'h000007b0344bc,
    48'h00000400597f8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b58,
    48'h00000400321e8,
    48'h0000040032288,
    48'h00000400ba2e4,
    48'h00000400ba2ec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032288,
    48'h00000400ba30c,
    48'h000007b0344b8,
    48'h00000400ba30c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0344b8,
    48'h000007b0337fc,
    48'h000007b0344b8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b034540,
    48'h000007b034380,
    48'h000004000e43c,
    48'h000007b034544,
    48'h000007b034544,
    48'h0000040059830,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b90,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6154,
    48'h00000400d615c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6174,
    48'h000007b0344b4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0344b4,
    48'h000007b034544,
    48'h000004005983c,
    48'h0000040059838,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b88,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b44,
    48'h00000400d5b4c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b64,
    48'h000007b034540,
    48'h00000400d5b64,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h00000400207cc,
    48'h000004002077c,
    48'h00000400207bc,
    48'h000007b0345fc,
    48'h000007b0345f8,
    48'h000007b0345f4,
    48'h000007b0345f0,
    48'h0000040020790,
    48'h00000400207cc,
    48'h000007b034380,
    48'h0000040020068,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h000007b034668,
    48'h000007b034380,
    48'h000004002048e,
    48'h000004000e43c,
    48'h000007b0345f4,
    48'h000007b034380,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f4,
    48'h0000040059838,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b4c,
    48'h000007b0345fc,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345fc,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h0000040059838,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b88,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b44,
    48'h00000400d5b4c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b64,
    48'h000007b0345f8,
    48'h00000400d5b64,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f8,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h0000040059770,
    48'h000007b0337fc,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h000007b034684,
    48'h0000040020054,
    48'h000007b034684,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0344b4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f4,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b0346bc,
    48'h000007b0344b4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h000007b0345f8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h000004007627c,
    48'h000007b0346bc,
    48'h000004007627c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0346bc,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0346b4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0344b4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b0344b4,
    48'h00000400f2ae0,
    48'h000007b0344b4,
    48'h00000400f2af8,
    48'h000007b0344b4,
    48'h00000400f2b00,
    48'h000007b0344b4,
    48'h00000400f2b0c,
    48'h000007b0344b4,
    48'h00000400f2b14,
    48'h000007b0344b4,
    48'h00000400f2b20,
    48'h000007b0344b4,
    48'h00000400f2b2c,
    48'h000007b0344b4,
    48'h00000400f2b38,
    48'h000007b0344b4,
    48'h00000400f2a20,
    48'h0000040020730,
    48'h000007b0344b4,
    48'h00000400f2a24,
    48'h000007b0344b4,
    48'h00000400f29f8,
    48'h000007b0344b4,
    48'h00000400f2aec,
    48'h000007b0344b4,
    48'h00000400f2a28,
    48'h000007b0344b4,
    48'h00000400f2a40,
    48'h000007b0344b4,
    48'h00000400f2a2c,
    48'h000007b0344b4,
    48'h00000400f2a34,
    48'h000007b0344b4,
    48'h00000400f2b44,
    48'h000007b0344b4,
    48'h00000400f2a4c,
    48'h000007b0344b4,
    48'h00000400f2a84,
    48'h000007b0337fc,
    48'h000007b0344b4,
    48'h0000040020068,
    48'h000007b0345f4,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03467c,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0347fc,
    48'h000007b0347f8,
    48'h000007b0347d4,
    48'h000007b0347d0,
    48'h0000040059780,
    48'h00000400f2a50,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761f0,
    48'h000007b0347d0,
    48'h00000400761f0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b0347d0,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040099500,
    48'h000007b0347f8,
    48'h0000040099500,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a4c,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034884,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h0000040020544,
    48'h000007b03490c,
    48'h000007b03490c,
    48'h000007b034984,
    48'h0000040020054,
    48'h000007b034984,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034884,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a4c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a4c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a4c,
    48'h000004003c00c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034884,
    48'h000007b0347d4,
    48'h000007b034884,
    48'h000007b034884,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a4c,
    48'h00000400323a4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b0348bc,
    48'h000007b0347d4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2a50,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761f0,
    48'h000007b0348bc,
    48'h00000400761f0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0348bc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0348b4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0347d4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347d4,
    48'h00000400f2b7c,
    48'h00000400f2b80,
    48'h00000400f2a4c,
    48'h0000040020468,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c00c,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c00c,
    48'h00000400f2b88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c74,
    48'h0000040045c74,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347f8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0347fc,
    48'h000007b0347f8,
    48'h000007b0347d4,
    48'h000007b0347d0,
    48'h0000040059780,
    48'h00000400f2a44,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076278,
    48'h000007b0347d0,
    48'h0000040076278,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b0347d0,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040099588,
    48'h000007b0347f8,
    48'h0000040099588,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a40,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034884,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h0000040020544,
    48'h000007b03490c,
    48'h000007b03490c,
    48'h000007b034984,
    48'h0000040020054,
    48'h000007b034984,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034884,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a40,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a40,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a40,
    48'h000004003c010,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034884,
    48'h000007b0347d4,
    48'h000007b034884,
    48'h000007b034884,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a40,
    48'h00000400323a8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b0348bc,
    48'h000007b0347d4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2a44,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076278,
    48'h000007b0348bc,
    48'h0000040076278,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0348bc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0348b4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0347d4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347d4,
    48'h00000400f3b84,
    48'h00000400f3b88,
    48'h00000400f2a40,
    48'h0000040020468,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c010,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c010,
    48'h00000400f3b90,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h0000040045c78,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347f8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h00000400f2a88,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0347fc,
    48'h000007b0347f8,
    48'h000007b0347d4,
    48'h000007b0347d0,
    48'h0000040059780,
    48'h00000400f2a88,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076274,
    48'h000007b0347d0,
    48'h0000040076274,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b0347d0,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040099584,
    48'h000007b0347f8,
    48'h0000040099584,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a84,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034884,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h0000040020544,
    48'h000007b03490c,
    48'h000007b03490c,
    48'h000007b034984,
    48'h0000040020054,
    48'h000007b034984,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034884,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a84,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a84,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a84,
    48'h000004003c014,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034884,
    48'h000007b0347d4,
    48'h000007b034884,
    48'h000007b034884,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a84,
    48'h00000400323ac,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b0348bc,
    48'h000007b0347d4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2a88,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076274,
    48'h000007b0348bc,
    48'h0000040076274,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0348bc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b03494c,
    48'h000007b034948,
    48'h000007b03494c,
    48'h000007b034948,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0348b4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0347d4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347d4,
    48'h00000400f3d0c,
    48'h00000400f3d10,
    48'h00000400f2a84,
    48'h0000040020468,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c014,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c014,
    48'h00000400f3d18,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c7c,
    48'h0000040045c7c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347f8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a84,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323ac,
    48'h00000400f2ab4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400f2a94,
    48'h000007b0337fc,
    48'h00000400f2a40,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b84,
    48'h000007b034724,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b88,
    48'h000007b034728,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b8c,
    48'h000007b03472c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b90,
    48'h000007b034730,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b94,
    48'h000007b034734,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b98,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h00000400f2a10,
    48'h00000400f2a5c,
    48'h000007b0337fc,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a28,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a28,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a28,
    48'h000004003c018,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a28,
    48'h00000400323b0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a28,
    48'h00000400323b0,
    48'h00000400f3e98,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a28,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3e94,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3ea8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3ea4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3e9c,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c018,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c80,
    48'h0000040045c80,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c80,
    48'h0000040045c80,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c80,
    48'h0000040045c80,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c80,
    48'h0000040045c80,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c80,
    48'h0000040045c80,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c80,
    48'h0000040045c80,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3e90,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3e94,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a28,
    48'h0000040045c80,
    48'h0000040045c80,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a28,
    48'h0000040045c80,
    48'h0000040045c80,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a28,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3e9c,
    48'h00000400f3e9c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3e98,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a2c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a2c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a2c,
    48'h000004003c01c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a2c,
    48'h00000400323b4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a2c,
    48'h00000400323b4,
    48'h00000400f4020,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a2c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f401c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f4030,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f402c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f4024,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c01c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c84,
    48'h0000040045c84,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c84,
    48'h0000040045c84,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c84,
    48'h0000040045c84,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c84,
    48'h0000040045c84,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c84,
    48'h0000040045c84,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c84,
    48'h0000040045c84,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f4018,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f401c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a2c,
    48'h0000040045c84,
    48'h0000040045c84,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a2c,
    48'h0000040045c84,
    48'h0000040045c84,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a2c,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f4024,
    48'h00000400f4024,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f4020,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347bc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b034838,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b034838,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b034944,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h0000040020544,
    48'h000007b0349cc,
    48'h000007b0349cc,
    48'h000007b034a44,
    48'h0000040020054,
    48'h000007b034a44,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034944,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a30,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a30,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a30,
    48'h000004003c020,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034944,
    48'h000007b034944,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a30,
    48'h00000400323b8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a30,
    48'h00000400323b8,
    48'h00000400f41a8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a30,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348c0,
    48'h000007b0348bc,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348c4,
    48'h000007b0348c0,
    48'h000007b0348bc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41a4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41b8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41b4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41ac,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c020,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c88,
    48'h0000040045c88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c88,
    48'h0000040045c88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c88,
    48'h0000040045c88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c88,
    48'h0000040045c88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c88,
    48'h0000040045c88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c88,
    48'h0000040045c88,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41a0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41a4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a30,
    48'h0000040045c88,
    48'h0000040045c88,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a30,
    48'h0000040045c88,
    48'h0000040045c88,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a30,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41ac,
    48'h00000400f41ac,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41a8,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a30,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h000007b0347bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a34,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a34,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a34,
    48'h000004003c024,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a34,
    48'h00000400323bc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a34,
    48'h00000400323bc,
    48'h00000400f4230,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a34,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f422c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f4240,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f423c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f4234,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c024,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c8c,
    48'h0000040045c8c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c8c,
    48'h0000040045c8c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c8c,
    48'h0000040045c8c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c8c,
    48'h0000040045c8c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c8c,
    48'h0000040045c8c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c8c,
    48'h0000040045c8c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f4228,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f422c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a34,
    48'h0000040045c8c,
    48'h0000040045c8c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a34,
    48'h0000040045c8c,
    48'h0000040045c8c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a34,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f4234,
    48'h00000400f4234,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f4230,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a34,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323bc,
    48'h00000400f2aa0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a38,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a38,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a38,
    48'h000004003c028,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a38,
    48'h00000400323c0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a38,
    48'h00000400323c0,
    48'h00000400f43b8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a38,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f43b4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f43c8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f43c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f43bc,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c028,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c90,
    48'h0000040045c90,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c90,
    48'h0000040045c90,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c90,
    48'h0000040045c90,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c90,
    48'h0000040045c90,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c90,
    48'h0000040045c90,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c90,
    48'h0000040045c90,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f43b0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f43b4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a38,
    48'h0000040045c90,
    48'h0000040045c90,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a38,
    48'h0000040045c90,
    48'h0000040045c90,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a38,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f43bc,
    48'h00000400f43bc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f43b8,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a38,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c0,
    48'h00000400f2aa4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034728,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a3c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a3c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a3c,
    48'h000004003c02c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a3c,
    48'h00000400323c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a3c,
    48'h00000400323c4,
    48'h00000400f4540,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a3c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f453c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f4550,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f454c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f4544,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c02c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c94,
    48'h0000040045c94,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c94,
    48'h0000040045c94,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c94,
    48'h0000040045c94,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c94,
    48'h0000040045c94,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c94,
    48'h0000040045c94,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c94,
    48'h0000040045c94,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f4538,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f453c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a3c,
    48'h0000040045c94,
    48'h0000040045c94,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a3c,
    48'h0000040045c94,
    48'h0000040045c94,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a3c,
    48'h000007b03472c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f4544,
    48'h00000400f4544,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f4540,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a3c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c4,
    48'h00000400f2aa8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a6c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a74,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a74,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a74,
    48'h000004003c030,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a74,
    48'h00000400323c8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a74,
    48'h00000400323c8,
    48'h00000400f46c8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a74,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f46c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f46d8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f46d4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f46cc,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c030,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c98,
    48'h0000040045c98,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c98,
    48'h0000040045c98,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c98,
    48'h0000040045c98,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c98,
    48'h0000040045c98,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c98,
    48'h0000040045c98,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c98,
    48'h0000040045c98,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f46c0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f46c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a74,
    48'h0000040045c98,
    48'h0000040045c98,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a74,
    48'h0000040045c98,
    48'h0000040045c98,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a74,
    48'h00000400f2a6c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f46cc,
    48'h00000400f46cc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f46c8,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a74,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323c8,
    48'h00000400f2aac,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a6c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0337fc,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347c4,
    48'h000007b0347c0,
    48'h000007b0347bc,
    48'h000007b0347b8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0348cc,
    48'h000007b0348cc,
    48'h0000040020544,
    48'h000007b03494c,
    48'h000007b03494c,
    48'h000007b0349c4,
    48'h0000040020054,
    48'h000007b0349c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2a78,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2a78,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2a78,
    48'h000004003c034,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0348c4,
    48'h000007b0348c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a78,
    48'h00000400323cc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2a78,
    48'h00000400323cc,
    48'h00000400f4750,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a78,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b034840,
    48'h000007b03483c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f474c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f4760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f475c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f4754,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c034,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c9c,
    48'h0000040045c9c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c9c,
    48'h0000040045c9c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c9c,
    48'h0000040045c9c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c9c,
    48'h0000040045c9c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c9c,
    48'h0000040045c9c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c9c,
    48'h0000040045c9c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f4748,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f474c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a78,
    48'h0000040045c9c,
    48'h0000040045c9c,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f2a78,
    48'h0000040045c9c,
    48'h0000040045c9c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a78,
    48'h00000400f2a6c,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f4754,
    48'h00000400f4754,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f4750,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a78,
    48'h000007b03474c,
    48'h000007b03474c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323cc,
    48'h00000400f2ab0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a60,
    48'h00000400f2a7c,
    48'h00000400f2a80,
    48'h00000400f2a70,
    48'h000007b0337fc,
    48'h00000400f2a5c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020344,
    48'h00000400f2a24,
    48'h000007b0337fc,
    48'h00000400f2ae4,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f2ae4,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761d8,
    48'h000007b034710,
    48'h00000400761d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994e8,
    48'h000007b034738,
    48'h00000400994e8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2ae0,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2ae0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2ae0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2ae0,
    48'h000004003c038,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2ae0,
    48'h00000400323d0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2ae4,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761d8,
    48'h000007b0347fc,
    48'h00000400761d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f47d4,
    48'h00000400f47d8,
    48'h00000400f2ae0,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c038,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c038,
    48'h00000400f47e0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca0,
    48'h0000040045ca0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f2afc,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761dc,
    48'h000007b034710,
    48'h00000400761dc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994ec,
    48'h000007b034738,
    48'h00000400994ec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2af8,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2af8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2af8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2af8,
    48'h000004003c03c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2af8,
    48'h00000400323d4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2afc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761dc,
    48'h000007b0347fc,
    48'h00000400761dc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f481c,
    48'h00000400f4820,
    48'h00000400f2af8,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c03c,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c03c,
    48'h00000400f4828,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca4,
    48'h0000040045ca4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f2b04,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761e0,
    48'h000007b034710,
    48'h00000400761e0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994f0,
    48'h000007b034738,
    48'h00000400994f0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2b00,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2b00,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2b00,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2b00,
    48'h000004003c040,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2b00,
    48'h00000400323d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2b04,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761e0,
    48'h000007b0347fc,
    48'h00000400761e0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f51a4,
    48'h00000400f51a8,
    48'h00000400f2b00,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c040,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c040,
    48'h00000400f51b0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ca8,
    48'h0000040045ca8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f2b10,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761e4,
    48'h000007b034710,
    48'h00000400761e4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994f4,
    48'h000007b034738,
    48'h00000400994f4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2b0c,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2b0c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2b0c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2b0c,
    48'h000004003c044,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2b0c,
    48'h00000400323dc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2b10,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761e4,
    48'h000007b0347fc,
    48'h00000400761e4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f5b2c,
    48'h00000400f5b30,
    48'h00000400f2b0c,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c044,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c044,
    48'h00000400f5b38,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cac,
    48'h0000040045cac,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f2b18,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761e8,
    48'h000007b034710,
    48'h00000400761e8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994f8,
    48'h000007b034738,
    48'h00000400994f8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2b14,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2b14,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2b14,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2b14,
    48'h000004003c048,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2b14,
    48'h00000400323e0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2b18,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761e8,
    48'h000007b0347fc,
    48'h00000400761e8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f5c74,
    48'h00000400f5c78,
    48'h00000400f2b14,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c048,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c048,
    48'h00000400f5c80,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb0,
    48'h0000040045cb0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f2b24,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761ec,
    48'h000007b034710,
    48'h00000400761ec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h00000400994fc,
    48'h000007b034738,
    48'h00000400994fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2b20,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f2b20,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f2b20,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f2b20,
    48'h000004003c04c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f2b20,
    48'h00000400323e4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f2b24,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761ec,
    48'h000007b0347fc,
    48'h00000400761ec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f5dbc,
    48'h00000400f5dc0,
    48'h00000400f2b20,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c04c,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c04c,
    48'h00000400f5dc8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb4,
    48'h0000040045cb4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h00000400f2b28,
    48'h000007b0337fc,
    48'h00000400f2b34,
    48'h000007b0337fc,
    48'h00000400f2b48,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f4,
    48'h0000040059830,
    48'h000007b0344b4,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03467c,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b0337fc,
    48'h000007b03467c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b90,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6154,
    48'h00000400d615c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03467c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6174,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000004002077c,
    48'h00000400207bc,
    48'h00000400207cc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034544,
    48'h0000040058f58,
    48'h0000040020344,
    48'h000007b0344b4,
    48'h00000400f2a24,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0344bc,
    48'h00000400597e8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b54,
    48'h00000400321e8,
    48'h0000040032284,
    48'h00000400a2b9c,
    48'h00000400a2ba4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032284,
    48'h00000400a2bc4,
    48'h000007b034404,
    48'h00000400a2bc4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0344b4,
    48'h00000400f2aec,
    48'h000007b034404,
    48'h00000400f2a10,
    48'h000007b0337fc,
    48'h000007b0344bc,
    48'h000007b0344b4,
    48'h000007b034404,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344c4,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344c4,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h00000400f2a5c,
    48'h00000400f2a10,
    48'h00000400f2a5c,
    48'h00000400f2a10,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b0345f8,
    48'h000007b0345f4,
    48'h000007b0345f0,
    48'h0000040020748,
    48'h000007b0345ec,
    48'h0000040058f58,
    48'h000007b0345ec,
    48'h000007b0345e8,
    48'h000007b034538,
    48'h00000400f2a28,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c80,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3e94,
    48'h00000400f3e9c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3eb0,
    48'h000007b03453c,
    48'h00000400f3eb0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03453c,
    48'h00000400f2a2c,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c84,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f401c,
    48'h00000400f4024,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f4038,
    48'h000007b0345f8,
    48'h00000400f4038,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345f8,
    48'h000007b0337fc,
    48'h00000400f2a40,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b84,
    48'h00000400f3b8c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3ba0,
    48'h000007b0345fc,
    48'h00000400f3ba0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0345fc,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b034600,
    48'h000007b034694,
    48'h000007b034690,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h0000040059770,
    48'h000007b034698,
    48'h0000040059774,
    48'h000007b03469c,
    48'h0000040059778,
    48'h000007b0346a0,
    48'h000004005977c,
    48'h000007b0346a4,
    48'h0000040059780,
    48'h000007b0346a8,
    48'h0000040059784,
    48'h000007b0346ac,
    48'h0000040059788,
    48'h000007b0346b0,
    48'h000004005978c,
    48'h000007b0346b4,
    48'h0000040059790,
    48'h000007b0346b8,
    48'h0000040059794,
    48'h000007b0346bc,
    48'h00000400f2a40,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b8c,
    48'h000007b034694,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034694,
    48'h00000400f2a40,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c78,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3b84,
    48'h00000400f3b8c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323a8,
    48'h00000400f3ba0,
    48'h000007b034690,
    48'h00000400f3ba0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346c4,
    48'h000007b03477c,
    48'h000007b034778,
    48'h000007b034754,
    48'h000007b034750,
    48'h000007b0346a8,
    48'h000007b034690,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761f4,
    48'h000007b034750,
    48'h00000400761f4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346b8,
    48'h000007b034750,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040099504,
    48'h000007b034778,
    48'h0000040099504,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03453c,
    48'h000007b034778,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034804,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03480c,
    48'h000007b03480c,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h000007b034904,
    48'h0000040020054,
    48'h000007b034904,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034804,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h000007b03453c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h000007b03453c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000007b03453c,
    48'h000004003c050,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034804,
    48'h000007b034754,
    48'h000007b034804,
    48'h000007b034804,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000007b03453c,
    48'h00000400323e8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034778,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03483c,
    48'h000007b034754,
    48'h000007b0337fc,
    48'h000007b0346a8,
    48'h000007b034690,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h00000400761f4,
    48'h000007b03483c,
    48'h00000400761f4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346b4,
    48'h000007b03483c,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b03484c,
    48'h000007b034848,
    48'h000007b034844,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h000007b0348cc,
    48'h000007b0348c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034834,
    48'h000007b0337fc,
    48'h000007b034698,
    48'h000007b034754,
    48'h000007b034698,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034754,
    48'h00000400f6144,
    48'h00000400f6148,
    48'h000007b03453c,
    48'h0000040020468,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c050,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c050,
    48'h00000400f6150,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cb8,
    48'h0000040045cb8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034778,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a20,
    48'h00000400f2a1c,
    48'h000007b0337fc,
    48'h00000400f2a28,
    48'h000007b03453c,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c80,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3e94,
    48'h00000400f3e9c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03473c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b0,
    48'h00000400f3eb0,
    48'h00000400f3eb0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a30,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41a8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c88,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41a4,
    48'h00000400f41ac,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b8,
    48'h00000400f41c0,
    48'h00000400f41c0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f2a2c,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b0346cc,
    48'h000007b0346c8,
    48'h000007b03473c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b0337fc,
    48'h000007b03473c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045c84,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f401c,
    48'h00000400f4024,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03473c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323b4,
    48'h00000400f4038,
    48'h00000400f4038,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400597c0,
    48'h00000400f29fc,
    48'h00000400f29f0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03453c,
    48'h000007b03460c,
    48'h000007b03460c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323e8,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020474,
    48'h0000040020474,
    48'h00000400f2a5c,
    48'h00000400f2a1c,
    48'h000007b0337fc,
    48'h00000400f29f0,
    48'h000007b03453c,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b0346c4,
    48'h000007b0346c0,
    48'h00000400207bc,
    48'h0000040020784,
    48'h000007b0346bc,
    48'h00000400205d8,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323e8,
    48'h000007b0346c0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346cc,
    48'h000007b0346cc,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323e8,
    48'h00000400f614c,
    48'h000007b0346c4,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0346c0,
    48'h000007b0346c4,
    48'h0000040020728,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h000007b0344b0,
    48'h000007b0337fc,
    48'h00000400207f8,
    48'h000007b0337fc,
    48'h0000040020788,
    48'h0000040020790,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0344b0,
    48'h000007b0344b4,
    48'h00000400f2a08,
    48'h000007b034384,
    48'h000007b0337fc,
    48'h000004002079c,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h00000400597e0,
    48'h000007b03437c,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03447c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032274,
    48'h00000400730c0,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b0337fc,
    48'h000007b03447c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b44,
    48'h00000400321e8,
    48'h0000040032274,
    48'h00000400730bc,
    48'h00000400730c4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032274,
    48'h00000400730d8,
    48'h00000400730d8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034400,
    48'h00000400597d0,
    48'h000007b03437c,
    48'h000007b034384,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03447c,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b034484,
    48'h000007b0337fc,
    48'h000007b03447c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b40,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b974,
    48'h000004005b97c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03447c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b99c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000004002079c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h00000400207d0,
    48'h00000400207bc,
    48'h00000400207cc,
    48'h000004002083c,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020090,
    48'h0000040020094,
    48'h0000040020078,
    48'h000004002007c,
    48'h0000040020080,
    48'h0000040020084,
    48'h0000040020088,
    48'h000004002008c,
    48'h000004002009c,
    48'h00000400200a0,
    48'h0000040020744,
    48'h000007b034298,
    48'h0000040020748,
    48'h000007b03429c,
    48'h000007b034294,
    48'h00000400207d0,
    48'h00000400207bc,
    48'h00000400207cc,
    48'h000004002083c,
    48'h000007b0342cc,
    48'h000007b0342c8,
    48'h000007b0342c4,
    48'h000007b0342c0,
    48'h000007b0342bc,
    48'h000007b0342b8,
    48'h000007b0342b4,
    48'h000007b0342b0,
    48'h000007b0342ac,
    48'h000007b0342a8,
    48'h000007b0342a4,
    48'h000007b0342a0,
    48'h000007b0342cc,
    48'h000007b0342c8,
    48'h000007b0342c4,
    48'h000007b0342c0,
    48'h000007b0342bc,
    48'h000007b0342b8,
    48'h000007b0342b4,
    48'h000007b0342b0,
    48'h000007b0342ac,
    48'h000007b0342a8,
    48'h000007b0342a4,
    48'h000007b0342a0,
    48'h000007b03438c,
    48'h000007b034388,
    48'h000007b034384,
    48'h000007b034380,
    48'h000007b03437c,
    48'h000007b034378,
    48'h000007b034374,
    48'h000007b034370,
    48'h000007b03436c,
    48'h000007b034368,
    48'h000007b034364,
    48'h000007b034360,
    48'h000007b03438c,
    48'h000007b034388,
    48'h000007b034384,
    48'h000007b034380,
    48'h000007b03437c,
    48'h000007b034378,
    48'h000007b034374,
    48'h000007b034370,
    48'h000007b03436c,
    48'h000007b034368,
    48'h000007b034364,
    48'h000007b034360,
    48'h00000400204ac,
    48'h00000400204b0,
    48'h00000400204b4,
    48'h00000400204b8,
    48'h00000400204bc,
    48'h00000400204c0,
    48'h00000400204c4,
    48'h00000400204c8,
    48'h00000400204cc,
    48'h00000400204d0,
    48'h00000400204d4,
    48'h00000400204d8,
    48'h00000400204dc,
    48'h00000400204e0,
    48'h00000400204e4,
    48'h00000400204e8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020438,
    48'h00000400f2970,
    48'h0000040020344,
    48'h0000040020360,
    48'h000004000e440,
    48'h00000400207cc,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000004002083c,
    48'h0000040020840,
    48'h000007b0337fc,
    48'h0000040020350,
    48'h000007b03429c,
    48'h000007b034298,
    48'h000007b0342cc,
    48'h000007b0342cc,
    48'h000007b034344,
    48'h000007b034340,
    48'h000007b03434c,
    48'h000007b03434c,
    48'h000007b0343c4,
    48'h000007b0343cc,
    48'h000007b0343cc,
    48'h000007b034428,
    48'h000007b03429c,
    48'h000004002048e,
    48'h000004000e43c,
    48'h000007b0343c4,
    48'h000007b03429c,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0343c4,
    48'h000007b034298,
    48'h000007b0343cc,
    48'h000007b0343c8,
    48'h000007b0343cc,
    48'h000007b0343c8,
    48'h000007b034294,
    48'h000007b0337fc,
    48'h00000400597d0,
    48'h000007b03444c,
    48'h000007b034448,
    48'h000007b03444c,
    48'h000007b034448,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h000007b0344cc,
    48'h000007b0344c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b40,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005b974,
    48'h000004005b97c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032270,
    48'h000004005bc70,
    48'h000007b034294,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034294,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03429c,
    48'h000004000e43c,
    48'h000007b034340,
    48'h000007b03434c,
    48'h000007b034348,
    48'h000007b03434c,
    48'h000007b034348,
    48'h000007b0343fc,
    48'h000007b0343f8,
    48'h000007b0343f4,
    48'h000007b0343f0,
    48'h000007b034298,
    48'h000007b03429c,
    48'h000004000e43c,
    48'h000007b0343fc,
    48'h000007b0343fc,
    48'h00000400597f8,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b03448c,
    48'h000007b034488,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b58,
    48'h00000400321e8,
    48'h0000040032288,
    48'h00000400ba2e4,
    48'h00000400ba2ec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032288,
    48'h00000400ba5e0,
    48'h000007b0343f8,
    48'h00000400ba5e0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0343f8,
    48'h000007b0337fc,
    48'h000007b0343f8,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b03440c,
    48'h000007b034408,
    48'h000007b034480,
    48'h000007b03429c,
    48'h000004000e43c,
    48'h000007b034484,
    48'h000007b034484,
    48'h0000040059830,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b03450c,
    48'h000007b034508,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b90,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d6154,
    48'h00000400d615c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322c0,
    48'h00000400d619c,
    48'h000007b0343f4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0343f4,
    48'h000007b034484,
    48'h000004005983c,
    48'h0000040059838,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b03450c,
    48'h000007b034508,
    48'h000007b03450c,
    48'h000007b034508,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b88,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b44,
    48'h00000400d5b4c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b8c,
    48'h000007b034480,
    48'h00000400d5b8c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03448c,
    48'h000007b034488,
    48'h000007b03448c,
    48'h000007b034488,
    48'h00000400207cc,
    48'h000004002077c,
    48'h00000400207bc,
    48'h000007b03453c,
    48'h000007b034538,
    48'h000007b034534,
    48'h000007b034530,
    48'h0000040020790,
    48'h00000400207cc,
    48'h000007b03429c,
    48'h0000040020068,
    48'h000007b03454c,
    48'h000007b03454c,
    48'h000007b0345a8,
    48'h000007b03429c,
    48'h000004002048e,
    48'h000004000e43c,
    48'h000007b034534,
    48'h000007b03429c,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034534,
    48'h0000040059838,
    48'h000007b03454c,
    48'h000007b03454c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b4c,
    48'h000007b03453c,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03453c,
    48'h000007b0337fc,
    48'h000007b034534,
    48'h0000040059838,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b88,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b44,
    48'h00000400d5b4c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400322b8,
    48'h00000400d5b8c,
    48'h000007b034538,
    48'h00000400d5b8c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034538,
    48'h000007b0337fc,
    48'h000007b034534,
    48'h0000040059770,
    48'h000007b0337fc,
    48'h000007b03454c,
    48'h000007b03454c,
    48'h000007b0345c4,
    48'h0000040020054,
    48'h000007b0345c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0343f4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034534,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b034540,
    48'h000007b0345fc,
    48'h000007b0343f4,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h000007b034538,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076434,
    48'h000007b0345fc,
    48'h0000040076434,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0345fc,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03460c,
    48'h000007b034608,
    48'h000007b034604,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0345f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b0343f4,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h000007b0343f4,
    48'h00000400f6738,
    48'h000007b0343f4,
    48'h00000400f6750,
    48'h000007b0343f4,
    48'h00000400f6758,
    48'h000007b0343f4,
    48'h00000400f6764,
    48'h000007b0343f4,
    48'h00000400f676c,
    48'h000007b0343f4,
    48'h00000400f6778,
    48'h000007b0343f4,
    48'h00000400f6784,
    48'h000007b0343f4,
    48'h00000400f6790,
    48'h000007b0343f4,
    48'h00000400f6678,
    48'h0000040020730,
    48'h000007b0343f4,
    48'h00000400f667c,
    48'h000007b0343f4,
    48'h00000400f6650,
    48'h000007b0343f4,
    48'h00000400f6744,
    48'h000007b0343f4,
    48'h00000400f6680,
    48'h000007b0343f4,
    48'h00000400f6698,
    48'h000007b0343f4,
    48'h00000400f6684,
    48'h000007b0343f4,
    48'h00000400f668c,
    48'h000007b0343f4,
    48'h00000400f679c,
    48'h000007b0343f4,
    48'h00000400f66a4,
    48'h000007b0343f4,
    48'h00000400f66dc,
    48'h000007b0337fc,
    48'h000007b0343f4,
    48'h0000040020068,
    48'h000007b034534,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b03454c,
    48'h000007b034548,
    48'h000007b034544,
    48'h000007b0345bc,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345c4,
    48'h000007b0345cc,
    48'h000007b0345c8,
    48'h000007b0345c4,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f66a8,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076424,
    48'h000007b034710,
    48'h0000040076424,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040099734,
    48'h000007b034738,
    48'h0000040099734,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f66a4,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f66a4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f66a4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f66a4,
    48'h000004003c054,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f66a4,
    48'h00000400323ec,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f66a8,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076424,
    48'h000007b0347fc,
    48'h0000040076424,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f67d4,
    48'h00000400f67d8,
    48'h00000400f66a4,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c054,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c054,
    48'h00000400f67e0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cbc,
    48'h0000040045cbc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f669c,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076430,
    48'h000007b034710,
    48'h0000040076430,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040099740,
    48'h000007b034738,
    48'h0000040099740,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f6698,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f6698,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f6698,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f6698,
    48'h000004003c058,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f6698,
    48'h00000400323f0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f669c,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040076430,
    48'h000007b0347fc,
    48'h0000040076430,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f77dc,
    48'h00000400f77e0,
    48'h00000400f6698,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c058,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c058,
    48'h00000400f77e8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc0,
    48'h0000040045cc0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020790,
    48'h000007b0337fc,
    48'h00000400f66e0,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b03473c,
    48'h000007b034738,
    48'h000007b034714,
    48'h000007b034710,
    48'h0000040059780,
    48'h00000400f66e0,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h000004007642c,
    48'h000007b034710,
    48'h000004007642c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040059790,
    48'h000007b034710,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h000007b0347cc,
    48'h000007b0347c8,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b50,
    48'h00000400321e8,
    48'h0000040032280,
    48'h0000040096fd4,
    48'h0000040096fdc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032280,
    48'h000004009973c,
    48'h000007b034738,
    48'h000004009973c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f66dc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b0347c4,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b0347cc,
    48'h000007b0347cc,
    48'h0000040020544,
    48'h000007b03484c,
    48'h000007b03484c,
    48'h000007b0348c4,
    48'h0000040020054,
    48'h000007b0348c4,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b0347c4,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f66dc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f66dc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f66dc,
    48'h000004003c05c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0347c4,
    48'h000007b034714,
    48'h000007b0347c4,
    48'h000007b0347c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f66dc,
    48'h00000400323f4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b034738,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b034744,
    48'h000007b034740,
    48'h000007b0347fc,
    48'h000007b034714,
    48'h000007b0337fc,
    48'h0000040059780,
    48'h00000400f66e0,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b48,
    48'h00000400321e8,
    48'h0000040032278,
    48'h0000040073cc4,
    48'h0000040073ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032278,
    48'h000004007642c,
    48'h000007b0347fc,
    48'h000004007642c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000004005978c,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b03488c,
    48'h000007b034888,
    48'h000007b03488c,
    48'h000007b034888,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045b4c,
    48'h00000400321e8,
    48'h000004003227c,
    48'h000004007f88c,
    48'h000004007f894,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h000004003227c,
    48'h00000400207bc,
    48'h0000040020784,
    48'h0000040020764,
    48'h0000040020820,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h000007b0347f4,
    48'h000007b0337fc,
    48'h0000040059770,
    48'h000007b034714,
    48'h0000040059770,
    48'h0000040020464,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034714,
    48'h00000400f7824,
    48'h00000400f7828,
    48'h00000400f66dc,
    48'h0000040020468,
    48'h000007b03474c,
    48'h000007b034748,
    48'h000007b03474c,
    48'h000007b034748,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c05c,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c05c,
    48'h00000400f7830,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc4,
    48'h0000040045cc4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034738,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f66dc,
    48'h000007b03468c,
    48'h000007b03468c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f4,
    48'h00000400f670c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400f66ec,
    48'h000007b0337fc,
    48'h00000400f6698,
    48'h000007b03468c,
    48'h000007b03468c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f0,
    48'h00000400f77dc,
    48'h000007b034664,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f0,
    48'h00000400f77e0,
    48'h000007b034668,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f0,
    48'h00000400f77e4,
    48'h000007b03466c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f0,
    48'h00000400f77e8,
    48'h000007b034670,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f0,
    48'h00000400f77ec,
    48'h000007b034674,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f0,
    48'h00000400f77f0,
    48'h000007b034678,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034668,
    48'h00000400f6668,
    48'h00000400f66b4,
    48'h000007b0337fc,
    48'h000007b034668,
    48'h000007b034678,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b034680,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b034680,
    48'h000007b0337fc,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b034704,
    48'h000007b034700,
    48'h000007b0346fc,
    48'h000007b0346f8,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b034704,
    48'h000007b034700,
    48'h000007b0346fc,
    48'h000007b0346f8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034804,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03480c,
    48'h000007b03480c,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h000007b034904,
    48'h0000040020054,
    48'h000007b034904,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034804,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f6680,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f6680,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f6680,
    48'h000004003c060,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034804,
    48'h000007b034804,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f6680,
    48'h00000400323f8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f6680,
    48'h00000400323f8,
    48'h00000400f7870,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f6680,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03477c,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03477c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f8,
    48'h00000400f786c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f8,
    48'h00000400f7880,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f8,
    48'h00000400f787c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f8,
    48'h00000400f7874,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c060,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc8,
    48'h0000040045cc8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc8,
    48'h0000040045cc8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc8,
    48'h0000040045cc8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc8,
    48'h0000040045cc8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc8,
    48'h0000040045cc8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cc8,
    48'h0000040045cc8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f8,
    48'h00000400f7868,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f8,
    48'h00000400f786c,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f6680,
    48'h0000040045cc8,
    48'h0000040045cc8,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f6680,
    48'h0000040045cc8,
    48'h0000040045cc8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f6680,
    48'h000007b03466c,
    48'h000007b03468c,
    48'h000007b03468c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f8,
    48'h00000400f7874,
    48'h00000400f7874,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323f8,
    48'h00000400f7870,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034668,
    48'h000007b034678,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b034680,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b034684,
    48'h000007b034680,
    48'h000007b0337fc,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b034704,
    48'h000007b034700,
    48'h000007b0346fc,
    48'h000007b0346f8,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b034704,
    48'h000007b034700,
    48'h000007b0346fc,
    48'h000007b0346f8,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034804,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03480c,
    48'h000007b03480c,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h000007b034904,
    48'h0000040020054,
    48'h000007b034904,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034804,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f6684,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f6684,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f6684,
    48'h000004003c064,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034804,
    48'h000007b034804,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f6684,
    48'h00000400323fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f6684,
    48'h00000400323fc,
    48'h00000400f78b8,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f6684,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03477c,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03477c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323fc,
    48'h00000400f78b4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323fc,
    48'h00000400f78c8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323fc,
    48'h00000400f78c4,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323fc,
    48'h00000400f78bc,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c064,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ccc,
    48'h0000040045ccc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ccc,
    48'h0000040045ccc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ccc,
    48'h0000040045ccc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ccc,
    48'h0000040045ccc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ccc,
    48'h0000040045ccc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045ccc,
    48'h0000040045ccc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323fc,
    48'h00000400f78b0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323fc,
    48'h00000400f78b4,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f6684,
    48'h0000040045ccc,
    48'h0000040045ccc,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f6684,
    48'h0000040045ccc,
    48'h0000040045ccc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f6684,
    48'h000007b03466c,
    48'h000007b03468c,
    48'h000007b03468c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323fc,
    48'h00000400f78bc,
    48'h00000400f78bc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400323fc,
    48'h00000400f78b8,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b03468c,
    48'h000007b034688,
    48'h000007b0346fc,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b034704,
    48'h000007b034700,
    48'h000007b03470c,
    48'h000007b034708,
    48'h000007b034704,
    48'h000007b034700,
    48'h000007b0337fc,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03477c,
    48'h000007b034778,
    48'h000007b03478c,
    48'h000007b034788,
    48'h000007b034784,
    48'h000007b034780,
    48'h000007b03477c,
    48'h000007b034778,
    48'h000007b0337fc,
    48'h000007b0337fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034884,
    48'h0000040020544,
    48'h0000040020764,
    48'h0000040020820,
    48'h0000040020544,
    48'h000007b03488c,
    48'h000007b03488c,
    48'h0000040020544,
    48'h000007b03490c,
    48'h000007b03490c,
    48'h000007b034984,
    48'h0000040020054,
    48'h000007b034984,
    48'h0000040020050,
    48'h0000040020014,
    48'h0000040020734,
    48'h0000040020004,
    48'h000004001fffc,
    48'h000004001ffe0,
    48'h000004001fffc,
    48'h000004002000c,
    48'h000004002000c,
    48'h0000040020014,
    48'h0000040020014,
    48'h0000040020018,
    48'h0000040020018,
    48'h000004002001c,
    48'h000004002001c,
    48'h0000040020058,
    48'h0000040020008,
    48'h00000400207e8,
    48'h00000400207bc,
    48'h000007b034884,
    48'h0000040020054,
    48'h000007b0337fc,
    48'h000004002004c,
    48'h000004002004c,
    48'h000004002076c,
    48'h0000040020774,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400207bc,
    48'h0000040020500,
    48'h000004003220c,
    48'h00000400f6688,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h000004003223c,
    48'h00000400f6688,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040020528,
    48'h0000040032250,
    48'h0000040032238,
    48'h0000040020528,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032250,
    48'h000004003223c,
    48'h000004003223c,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032254,
    48'h000004003bea4,
    48'h000004003bea4,
    48'h000004002052c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032258,
    48'h0000040045b0c,
    48'h0000040045b0c,
    48'h000004002052c,
    48'h0000040020530,
    48'h0000040020530,
    48'h0000040020534,
    48'h0000040020534,
    48'h0000040020500,
    48'h00000400321ec,
    48'h00000400f6688,
    48'h000004003c068,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b034884,
    48'h000007b034884,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f6688,
    48'h0000040032400,
    48'h0000040020500,
    48'h00000400321e8,
    48'h00000400f6688,
    48'h0000040032400,
    48'h00000400f7900,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f6688,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b0347fc,
    48'h000007b03480c,
    48'h000007b034808,
    48'h000007b034804,
    48'h000007b034800,
    48'h000007b0347fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h00000400f78fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h00000400f7910,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h00000400f790c,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h00000400f7904,
    48'h0000040020500,
    48'h00000400321ec,
    48'h000004003c068,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cd0,
    48'h0000040045cd0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cd0,
    48'h0000040045cd0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cd0,
    48'h0000040045cd0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cd0,
    48'h0000040045cd0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cd0,
    48'h0000040045cd0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h0000040045cd0,
    48'h0000040045cd0,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h00000400f78f8,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h00000400f78fc,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h000007b0337fc,
    48'h00000400207bc,
    48'h0000040020550,
    48'h0000040020784,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f6688,
    48'h0000040045cd0,
    48'h0000040045cd0,
    48'h0000040020500,
    48'h00000400321f0,
    48'h00000400f6688,
    48'h0000040045cd0,
    48'h0000040045cd0,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f6688,
    48'h000007b03470c,
    48'h000007b03470c,
    48'h0000040020504,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h00000400f7904,
    48'h00000400f7904,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h00000400f7900,
    48'h000007b0337fc,
    48'h0000040020508,
    48'h000007b0337fc,
    48'h0000040020760,
    48'h0000040020760,
    48'h00000400f6688,
    48'h000007b03470c,
    48'h000007b03470c,
    48'h0000040020530,
    48'h0000040020504,
    48'h000007b0337fc,
    48'h0000040020500,
    48'h00000400321e8,
    48'h0000040032400,
    48'h000007b0346fc
    };
endmodule