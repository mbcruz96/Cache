
parameter SIZE = 20000;
module trace_addr(
    reg[47:0] test_addrs[0:SIZE-1]);
    
    assign test_addrs = 
    {
    48'h00000400341a0,
    48'h0000000dfcfa8,
    48'h000007b034dd4,
    48'h0000000df7c48,
    48'h000007b034dd4,
    48'h00000423aebbc,
    48'h00000423aebb8,
    48'h00000423aebbc,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423aeb9c,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423aeba0,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df8a70,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9f10,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8a74,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000df9f14,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h00000423aeb90,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000040139dd0,
    48'h00000423aeb92,
    48'h00000423aeb94,
    48'h00000423aeb88,
    48'h00000423aeb88,
    48'h00000423aeb88,
    48'h00000423aeb88,
    48'h00000423aeb8c,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h00000423aeb88,
    48'h0000040022e80,
    48'h00000423aeb88,
    48'h000004214c9d4,
    48'h0000040002178,
    48'h0000000384130,
    48'h00000423aeb8c,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h00000401367d0,
    48'h000007b0345e4,
    48'h00000423aeb8c,
    48'h00000423aeb94,
    48'h0000040022e80,
    48'h0000040139dd0,
    48'h00000423aeb9c,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000004013893c,
    48'h00000423aeb80,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423aeb82,
    48'h00000423aeb84,
    48'h00000423aeb70,
    48'h00000423aeb70,
    48'h00000423aeb70,
    48'h00000423aeb70,
    48'h00000423aeb70,
    48'h00000423aeb74,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423aeb78,
    48'h00000423aeb68,
    48'h00000423aeb6c,
    48'h00000423aeb70,
    48'h00000423aeb78,
    48'h00000423aeb68,
    48'h00000423aeb74,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h00000423aeba0,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h00000423aeb90,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b034d58,
    48'h0000000df84d5,
    48'h000007b034dfc,
    48'h00000423aeb90,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h00000423aeb90,
    48'h0000000df84d6,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h00000423aeb80,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034c9c,
    48'h0000040139a84,
    48'h000007b034c9c,
    48'h00000423aeb80,
    48'h0000000df84e5,
    48'h000007b034c9c,
    48'h0000040139bac,
    48'h000007b034c9c,
    48'h00000423aeb80,
    48'h0000000df84e6,
    48'h000007b034c9c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034c9c,
    48'h00000423aeb80,
    48'h0000000df84e7,
    48'h000007b034dfc,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h0000000df84e8,
    48'h00000423aeb80,
    48'h0000000df84e9,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h0000000df84ea,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423aeb9c,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423aeba0,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h00000423aeb90,
    48'h00000423aeb90,
    48'h00000423aeb90,
    48'h000007b034ce0,
    48'h000007b034d58,
    48'h00000423aeba8,
    48'h000007b034d58,
    48'h000007b034d58,
    48'h0000040138938,
    48'h000007b034ce0,
    48'h000007b034e94,
    48'h000007b034d58,
    48'h000007b034e90,
    48'h000007b034d58,
    48'h000007b034da8,
    48'h000007b034e8c,
    48'h000007b034dcc,
    48'h0000000dfb1df,
    48'h000007b034e88,
    48'h000007b034e84,
    48'h0000040139dd0,
    48'h000007b034e90,
    48'h000007b034e8c,
    48'h000007b034e88,
    48'h000007b034e94,
    48'h00000423aeb90,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423aeb9c,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000040022cb0,
    48'h0000040022e88,
    48'h000007b034cf8,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h000007b034ce4,
    48'h000007b034d5c,
    48'h000007b034d5c,
    48'h000004013893c,
    48'h000007b034d5c,
    48'h000007b034ce4,
    48'h000007b034e94,
    48'h000007b034d5c,
    48'h000007b034dac,
    48'h000007b034e90,
    48'h000007b034d5c,
    48'h000007b034e8c,
    48'h000007b034dcc,
    48'h0000000dfb1e0,
    48'h000007b034e88,
    48'h000007b034e84,
    48'h0000040139dd4,
    48'h000007b034e90,
    48'h000007b034e8c,
    48'h000007b034e88,
    48'h000007b034e94,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb82,
    48'h0000040136800,
    48'h0000040139540,
    48'h000004214c780,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040139540,
    48'h000004214c780,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c494,
    48'h000004214c69c,
    48'h0000040139544,
    48'h000004214c344,
    48'h000004013885c,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136514,
    48'h000004214c781,
    48'h000004214c599,
    48'h00000423aeba0,
    48'h0000040136800,
    48'h0000040138f44,
    48'h00000423aeba0,
    48'h0000040022cb0,
    48'h000007b034cfc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000004214c69c,
    48'h0000040136800,
    48'h0000040138eb0,
    48'h000007b034dcc,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000007b03451c,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423aebaa,
    48'h000007b034390,
    48'h000007b0344a8,
    48'h000007b034400,
    48'h000007b0344e0,
    48'h000007b034394,
    48'h000007b0344ac,
    48'h000007b034404,
    48'h000007b0344e4,
    48'h000007b034398,
    48'h000007b0344b0,
    48'h000007b034408,
    48'h000007b0344e8,
    48'h000007b03439c,
    48'h000007b0344b4,
    48'h000007b03440c,
    48'h000007b0344ec,
    48'h000007b0343a0,
    48'h000007b0344b8,
    48'h000007b034410,
    48'h000007b0344f0,
    48'h000007b0343a4,
    48'h000007b0344bc,
    48'h000007b034414,
    48'h000007b0344f4,
    48'h000007b0343a8,
    48'h000007b0344c0,
    48'h000007b034418,
    48'h000007b0344f8,
    48'h000007b0343ac,
    48'h000007b0344c4,
    48'h000007b03441c,
    48'h000007b0344fc,
    48'h000007b0343b0,
    48'h000007b0344c8,
    48'h000007b034420,
    48'h000007b034500,
    48'h000007b0343b4,
    48'h000007b0344cc,
    48'h000007b034424,
    48'h000007b034504,
    48'h000007b0343b8,
    48'h000007b0344d0,
    48'h000007b034428,
    48'h000007b034508,
    48'h000007b0343bc,
    48'h000007b0344d4,
    48'h000007b03442c,
    48'h000007b03450c,
    48'h000007b0343c0,
    48'h000007b0344d8,
    48'h000007b034430,
    48'h000007b034510,
    48'h000007b0343c4,
    48'h000007b0344dc,
    48'h000007b034434,
    48'h000007b034514,
    48'h00000423aebb4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423aebe0,
    48'h00000423aebe0,
    48'h00000423aebec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423aec30,
    48'h00000423aec30,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423aec40,
    48'h00000423aec20,
    48'h000004214c8a8,
    48'h00000423aec44,
    48'h00000423aec44,
    48'h000007b034dcc,
    48'h0000000dfd2f8,
    48'h000007b034dd4,
    48'h0000000df7f98,
    48'h000007b034dd4,
    48'h00000423aec44,
    48'h00000423aec40,
    48'h00000423aec44,
    48'h0000040002984,
    48'h0000040139dd0,
    48'h00000423aec24,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423aec28,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df9b00,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000dfafa0,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df9b04,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000dfafa4,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df8778,
    48'h0000000df8779,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84f8,
    48'h0000000df84f9,
    48'h0000040138938,
    48'h00000423aec18,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df8778,
    48'h0000040138938,
    48'h0000040139dd0,
    48'h00000423aec1a,
    48'h00000423aec1c,
    48'h000004239fdc8,
    48'h000004239fdc8,
    48'h000004239fdc8,
    48'h0000040022e80,
    48'h000004239fdc8,
    48'h00000423aec1c,
    48'h0000040022e80,
    48'h0000040139dd0,
    48'h00000423aec24,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000004013893c,
    48'h00000423aec10,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84f8,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h00000423aec18,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df8778,
    48'h0000000df8778,
    48'h000007b034dfc,
    48'h00000423aec18,
    48'h00000423aec18,
    48'h00000423aec1a,
    48'h00000423aec1c,
    48'h000007b034f50,
    48'h000004239fdc8,
    48'h000004239fdc8,
    48'h00000423aec18,
    48'h00000423aec18,
    48'h000007b034df4,
    48'h0000000df8779,
    48'h000007b034c68,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h00000423aec10,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84f8,
    48'h0000000df84f8,
    48'h000007b034dfc,
    48'h00000423aec10,
    48'h000007b034c9c,
    48'h0000040139a98,
    48'h000007b034c9c,
    48'h00000423aec10,
    48'h0000000df84f9,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423aec24,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423aec28,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h00000423aec18,
    48'h00000423aec18,
    48'h00000423aec18,
    48'h000007b034ce0,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423aec10,
    48'h00000423aec10,
    48'h00000423aec10,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df83b8,
    48'h0000040136800,
    48'h00000423aec3c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423aec78,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423aec88,
    48'h00000423aec68,
    48'h00000423aec6c,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h00000423aec70,
    48'h00000423aec58,
    48'h00000423aec68,
    48'h00000423aec68,
    48'h00000423aec70,
    48'h00000423aec58,
    48'h00000423aec68,
    48'h000004214c8a8,
    48'h00000423aec8c,
    48'h00000423aec8c,
    48'h000007b034dcc,
    48'h0000000dfd064,
    48'h000007b034dd4,
    48'h0000000df7d04,
    48'h000007b034dd4,
    48'h00000423aec8c,
    48'h00000423aec88,
    48'h00000423aec8c,
    48'h00000400026f0,
    48'h0000040139dd0,
    48'h00000423aec6c,
    48'h0000040138938,
    48'h00000423aec70,
    48'h0000040139dd4,
    48'h00000423aec5c,
    48'h000004013893c,
    48'h00000423aec70,
    48'h0000040139dd8,
    48'h00000423aec60,
    48'h0000040138940,
    48'h000007b034dcc,
    48'h0000000df8e1c,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000dfa2bc,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8e20,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000dfa2c0,
    48'h000007b034dac,
    48'h000007b034dcc,
    48'h0000000df8e24,
    48'h000007b034c58,
    48'h000007b034c70,
    48'h0000000dfa2c4,
    48'h000007b034db0,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df863c,
    48'h0000000df863d,
    48'h0000000df863e,
    48'h0000000df863f,
    48'h0000000df8640,
    48'h0000000df8641,
    48'h0000000df8642,
    48'h0000000df8643,
    48'h0000000df8644,
    48'h0000000df8645,
    48'h0000000df8646,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df8648,
    48'h0000000df8649,
    48'h0000040138938,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034d71,
    48'h0000040138938,
    48'h0000040138940,
    48'h0000042351e38,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h000007b034d72,
    48'h0000000df864a,
    48'h0000000df864b,
    48'h0000040138938,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034d71,
    48'h0000040138938,
    48'h0000040138940,
    48'h0000042351e38,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h000007b034d72,
    48'h0000000df864c,
    48'h0000000df864d,
    48'h0000000df864e,
    48'h0000000df864f,
    48'h0000000df8650,
    48'h0000000df8651,
    48'h0000000df8652,
    48'h0000040138940,
    48'h000007b034d98,
    48'h000007b034c70,
    48'h0000000df8654,
    48'h0000000df8655,
    48'h0000000df8656,
    48'h0000000df8657,
    48'h0000000df8658,
    48'h0000000df8659,
    48'h0000000df865a,
    48'h0000000df865b,
    48'h0000000df865c,
    48'h0000000df865d,
    48'h0000000df865e,
    48'h0000000df865f,
    48'h0000000df8660,
    48'h0000000df8661,
    48'h0000000df8662,
    48'h0000000df8663,
    48'h0000000df8664,
    48'h0000000df8665,
    48'h0000000df8666,
    48'h0000040138938,
    48'h0000042351e38,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df863c,
    48'h0000040138938,
    48'h0000042351e3c,
    48'h00000401367d0,
    48'h000007b0345e4,
    48'h0000040136428,
    48'h000007b034a64,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df8648,
    48'h000004013893c,
    48'h0000042351e3c,
    48'h00000401367d0,
    48'h000007b0345e4,
    48'h0000040136428,
    48'h000007b034a64,
    48'h0000040138940,
    48'h00000423aec50,
    48'h000007b034d60,
    48'h000007b034c88,
    48'h000007b034c70,
    48'h0000000df8654,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042351e38,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df863c,
    48'h0000000df863c,
    48'h000007b034d58,
    48'h0000000df863d,
    48'h000007b034dfc,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h0000042351e38,
    48'h0000042351e38,
    48'h0000000df863e,
    48'h000007b034c68,
    48'h000007b034cc0,
    48'h000007b034cb8,
    48'h000007b034de4,
    48'h0000042351e38,
    48'h000007b034c98,
    48'h000007b034cc8,
    48'h000007b034de4,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df8648,
    48'h0000000df8648,
    48'h0000000df8649,
    48'h000007b034ccc,
    48'h000007b034ddc,
    48'h000007b034d71,
    48'h000007b034cb0,
    48'h000007b034c98,
    48'h000007b034c9c,
    48'h0000000df864a,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034cb9,
    48'h0000042351e38,
    48'h000007b034c9c,
    48'h000007b034ccc,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h00000423aec50,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df8654,
    48'h0000000df8654,
    48'h000007b034ca0,
    48'h0000040139a84,
    48'h000007b034ca0,
    48'h00000423aec50,
    48'h0000000df8655,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8656,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8657,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8658,
    48'h00000423aec50,
    48'h0000000df8659,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034cba,
    48'h00000423aec50,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034dec,
    48'h000007b034de4,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042351e38,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df863f,
    48'h0000000df863f,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042351e38,
    48'h0000040138938,
    48'h0000042351e3a,
    48'h000007b034c98,
    48'h0000042351e3c,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df8640,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df864b,
    48'h0000000df864b,
    48'h000007b034ccc,
    48'h000007b034ddc,
    48'h000007b034d71,
    48'h000007b034cb0,
    48'h000007b034c98,
    48'h000007b034c9c,
    48'h0000000df864c,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h00000423aec50,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df865a,
    48'h0000000df865a,
    48'h000007b034dfc,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h0000000df865b,
    48'h000007b034ca0,
    48'h0000040139a98,
    48'h000007b034ca0,
    48'h00000423aec50,
    48'h0000000df865c,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df865d,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df865e,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df865f,
    48'h00000423aec50,
    48'h0000000df8660,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034cba,
    48'h00000423aec50,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034dec,
    48'h000007b034de4,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb0,
    48'h000007b034d40,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb1,
    48'h000007b034d41,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ca0,
    48'h000007b034ce8,
    48'h000007b034cb2,
    48'h000007b034d42,
    48'h000007b034cba,
    48'h000007b034d4a,
    48'h000007b034cd0,
    48'h000007b034d18,
    48'h000007b034cc2,
    48'h000007b034d52,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042351e38,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df8641,
    48'h0000000df8641,
    48'h000007b034dec,
    48'h0000000df8642,
    48'h000007b034c98,
    48'h0000040139a94,
    48'h000007b034c98,
    48'h0000042351e38,
    48'h0000040138938,
    48'h0000042351e3a,
    48'h000007b034c98,
    48'h0000042351e3c,
    48'h00000400024b0,
    48'h0000040001fac,
    48'h0000000df8643,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df864d,
    48'h0000000df864d,
    48'h000007b034c9c,
    48'h0000040139a94,
    48'h000007b034c9c,
    48'h0000042351e38,
    48'h000004013893c,
    48'h0000042351e3a,
    48'h000007b034c9c,
    48'h0000042351e3c,
    48'h00000400024b0,
    48'h0000040001fac,
    48'h0000000df864e,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h00000423aec50,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df8661,
    48'h0000000df8661,
    48'h000007b034ca0,
    48'h0000040139a98,
    48'h000007b034ca0,
    48'h00000423aec50,
    48'h0000000df8662,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8663,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8664,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034dfc,
    48'h000007b034cb2,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034d94,
    48'h000004013893c,
    48'h000007b034d98,
    48'h0000040138940,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034d42,
    48'h000007b034ca0,
    48'h000007b034ce8,
    48'h000007b034cba,
    48'h000007b034d4a,
    48'h000007b034cd0,
    48'h000007b034d18,
    48'h000007b034cc2,
    48'h000007b034d52,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d30,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d42,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423aec6c,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423aec5c,
    48'h000007b034cfc,
    48'h0000040139dd8,
    48'h000007b034d98,
    48'h00000423aec60,
    48'h000007b034d00,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d42,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042351e38,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h0000042351e38,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042351e38,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h0000042351e38,
    48'h000007b034d42,
    48'h000007b034d30,
    48'h000007b034d18,
    48'h00000400015a4,
    48'h0000040138940,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8124,
    48'h0000040136800,
    48'h00000423aec84,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423afca8,
    48'h00000423afca8,
    48'h00000423afcb4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423ae400,
    48'h00000423ae400,
    48'h00000423ae40c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423afcf8,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afd08,
    48'h00000423afce8,
    48'h00000423afcec,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423afcf0,
    48'h00000423afce0,
    48'h00000423afce8,
    48'h00000423afce8,
    48'h00000423afcf0,
    48'h00000423afce0,
    48'h00000423afce8,
    48'h000004214c8a8,
    48'h00000423afd0c,
    48'h00000423afd0c,
    48'h000007b034dcc,
    48'h0000000dfcfa8,
    48'h000007b034dd4,
    48'h0000000df7c48,
    48'h000007b034dd4,
    48'h00000423afd0c,
    48'h00000423afd08,
    48'h00000423afd0c,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423afcec,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423afcf0,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df8a70,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9f10,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8a74,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000df9f14,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040136428,
    48'h000007b034a50,
    48'h000004013893c,
    48'h00000423afce0,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423afce2,
    48'h00000423afce4,
    48'h00000423afcd0,
    48'h00000423afcd0,
    48'h00000423afcd0,
    48'h00000423afcd0,
    48'h00000423afcd0,
    48'h00000423afcd4,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423afcd8,
    48'h00000423afcc8,
    48'h00000423afccc,
    48'h00000423afcd0,
    48'h00000423afcd8,
    48'h00000423afcc8,
    48'h00000423afcd4,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h00000423afcf0,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b034d58,
    48'h0000000df84d5,
    48'h000007b034dfc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354d90,
    48'h0000040138938,
    48'h0000042354d92,
    48'h000007b034c98,
    48'h0000042354d94,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h00000423afce0,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034c9c,
    48'h0000040139a84,
    48'h000007b034c9c,
    48'h00000423afce0,
    48'h0000000df84e5,
    48'h000007b034c9c,
    48'h0000040139bac,
    48'h000007b034c9c,
    48'h00000423afce0,
    48'h0000000df84e6,
    48'h000007b034c9c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034c9c,
    48'h00000423afce0,
    48'h0000000df84e7,
    48'h000007b034dfc,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h0000000df84e8,
    48'h00000423afce0,
    48'h0000000df84e9,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h0000000df84ea,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423afcec,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423afcf0,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d90,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h000007b034ce4,
    48'h000007b034d5c,
    48'h000007b034d5c,
    48'h000004013893c,
    48'h000007b034d5c,
    48'h000007b034ce4,
    48'h000007b034e94,
    48'h000007b034d5c,
    48'h000007b034dac,
    48'h000007b034e90,
    48'h000007b034d5c,
    48'h000007b034e8c,
    48'h000007b034dcc,
    48'h0000000dfb1e0,
    48'h000007b034e88,
    48'h000007b034e84,
    48'h0000040139dd4,
    48'h000007b034e90,
    48'h000007b034e8c,
    48'h000007b034e88,
    48'h000007b034e94,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423afcf0,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423afcf0,
    48'h0000040022cb0,
    48'h000007b034cfc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000007b03451c,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423afcfa,
    48'h000007b034390,
    48'h000007b0344a8,
    48'h000007b034400,
    48'h000007b0344e0,
    48'h000007b034394,
    48'h000007b0344ac,
    48'h000007b034404,
    48'h000007b0344e4,
    48'h000007b034398,
    48'h000007b0344b0,
    48'h000007b034408,
    48'h000007b0344e8,
    48'h000007b03439c,
    48'h000007b0344b4,
    48'h000007b03440c,
    48'h000007b0344ec,
    48'h000007b0343a0,
    48'h000007b0344b8,
    48'h000007b034410,
    48'h000007b0344f0,
    48'h000007b0343a4,
    48'h000007b0344bc,
    48'h000007b034414,
    48'h000007b0344f4,
    48'h000007b0343a8,
    48'h000007b0344c0,
    48'h000007b034418,
    48'h000007b0344f8,
    48'h000007b0343ac,
    48'h000007b0344c4,
    48'h000007b03441c,
    48'h000007b0344fc,
    48'h000007b0343b0,
    48'h000007b0344c8,
    48'h000007b034420,
    48'h000007b034500,
    48'h000007b0343b4,
    48'h000007b0344cc,
    48'h000007b034424,
    48'h000007b034504,
    48'h000007b0343b8,
    48'h000007b0344d0,
    48'h000007b034428,
    48'h000007b034508,
    48'h000007b0343bc,
    48'h000007b0344d4,
    48'h000007b03442c,
    48'h000007b03450c,
    48'h000007b0343c0,
    48'h000007b0344d8,
    48'h000007b034430,
    48'h000007b034510,
    48'h000007b0343c4,
    48'h000007b0344dc,
    48'h000007b034434,
    48'h000007b034514,
    48'h00000423afd04,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423afd50,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afd60,
    48'h00000423afd40,
    48'h00000423afd44,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000423afd48,
    48'h00000423afd38,
    48'h00000423afd40,
    48'h00000423afd40,
    48'h00000423afd48,
    48'h00000423afd38,
    48'h00000423afd40,
    48'h000004214c8a8,
    48'h00000423afd64,
    48'h00000423afd64,
    48'h000007b034dcc,
    48'h0000000dfcfa8,
    48'h000007b034dd4,
    48'h0000000df7c48,
    48'h000007b034dd4,
    48'h00000423afd64,
    48'h00000423afd60,
    48'h00000423afd64,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423afd44,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423afd48,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df8a70,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9f10,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8a74,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000df9f14,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354d00,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040136428,
    48'h000007b034a54,
    48'h000004013893c,
    48'h00000423afd38,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423afd3a,
    48'h00000423afd3c,
    48'h00000423afd28,
    48'h00000423afd28,
    48'h00000423afd28,
    48'h00000423afd28,
    48'h00000423afd28,
    48'h00000423afd2c,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000423afd30,
    48'h00000423afd20,
    48'h00000423afd24,
    48'h00000423afd28,
    48'h00000423afd30,
    48'h00000423afd20,
    48'h00000423afd2c,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040139dd4,
    48'h00000423afd48,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354d00,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b034d58,
    48'h0000000df84d5,
    48'h000007b034dfc,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354d00,
    48'h0000040138938,
    48'h0000042354d02,
    48'h000007b034c98,
    48'h0000042354d04,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h00000423afd38,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034c9c,
    48'h0000040139a84,
    48'h000007b034c9c,
    48'h00000423afd38,
    48'h0000000df84e5,
    48'h000007b034c9c,
    48'h0000040139bac,
    48'h000007b034c9c,
    48'h00000423afd38,
    48'h0000000df84e6,
    48'h000007b034c9c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034c9c,
    48'h00000423afd38,
    48'h0000000df84e7,
    48'h000007b034dfc,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h0000000df84e8,
    48'h00000423afd38,
    48'h0000000df84e9,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h0000000df84ea,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423afd44,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423afd48,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042354d00,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h000007b034ce4,
    48'h000007b034d5c,
    48'h000007b034d5c,
    48'h000004013893c,
    48'h000007b034d5c,
    48'h000007b034ce4,
    48'h000007b034e94,
    48'h000007b034d5c,
    48'h000007b034dac,
    48'h000007b034e90,
    48'h000007b034d5c,
    48'h000007b034e8c,
    48'h000007b034dcc,
    48'h0000000dfb1e0,
    48'h000007b034e88,
    48'h000007b034e84,
    48'h0000040139dd4,
    48'h000007b034e90,
    48'h000007b034e8c,
    48'h000007b034e88,
    48'h000007b034e94,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd3a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423afd48,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423afd48,
    48'h0000040022cb0,
    48'h000007b034cfc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000007b03451c,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423afd52,
    48'h000007b034390,
    48'h000007b0344a8,
    48'h000007b034400,
    48'h000007b0344e0,
    48'h000007b034394,
    48'h000007b0344ac,
    48'h000007b034404,
    48'h000007b0344e4,
    48'h000007b034398,
    48'h000007b0344b0,
    48'h000007b034408,
    48'h000007b0344e8,
    48'h000007b03439c,
    48'h000007b0344b4,
    48'h000007b03440c,
    48'h000007b0344ec,
    48'h000007b0343a0,
    48'h000007b0344b8,
    48'h000007b034410,
    48'h000007b0344f0,
    48'h000007b0343a4,
    48'h000007b0344bc,
    48'h000007b034414,
    48'h000007b0344f4,
    48'h000007b0343a8,
    48'h000007b0344c0,
    48'h000007b034418,
    48'h000007b0344f8,
    48'h000007b0343ac,
    48'h000007b0344c4,
    48'h000007b03441c,
    48'h000007b0344fc,
    48'h000007b0343b0,
    48'h000007b0344c8,
    48'h000007b034420,
    48'h000007b034500,
    48'h000007b0343b4,
    48'h000007b0344cc,
    48'h000007b034424,
    48'h000007b034504,
    48'h000007b0343b8,
    48'h000007b0344d0,
    48'h000007b034428,
    48'h000007b034508,
    48'h000007b0343bc,
    48'h000007b0344d4,
    48'h000007b03442c,
    48'h000007b03450c,
    48'h000007b0343c0,
    48'h000007b0344d8,
    48'h000007b034430,
    48'h000007b034510,
    48'h000007b0343c4,
    48'h000007b0344dc,
    48'h000007b034434,
    48'h000007b034514,
    48'h00000423afd5c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423afda8,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afdb8,
    48'h00000423afd80,
    48'h00000423afd84,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423afd88,
    48'h00000423afd70,
    48'h00000423afd80,
    48'h00000423afd80,
    48'h00000423afd88,
    48'h00000423afd70,
    48'h00000423afd80,
    48'h000004214c8a8,
    48'h00000423afdbc,
    48'h00000423afdbc,
    48'h000007b034dcc,
    48'h0000000dfd064,
    48'h000007b034dd4,
    48'h0000000df7d04,
    48'h000007b034dd4,
    48'h00000423afdbc,
    48'h00000423afdb8,
    48'h00000423afdbc,
    48'h00000400026f0,
    48'h0000040139dd0,
    48'h00000423afd84,
    48'h0000040138938,
    48'h00000423afd88,
    48'h0000040139dd4,
    48'h00000423afd74,
    48'h000004013893c,
    48'h00000423afd88,
    48'h0000040139dd8,
    48'h00000423afd78,
    48'h0000040138940,
    48'h000007b034dcc,
    48'h0000000df8e1c,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000dfa2bc,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8e20,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000dfa2c0,
    48'h000007b034dac,
    48'h000007b034dcc,
    48'h0000000df8e24,
    48'h000007b034c58,
    48'h000007b034c70,
    48'h0000000dfa2c4,
    48'h000007b034db0,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df863c,
    48'h0000000df863d,
    48'h0000000df863e,
    48'h0000000df863f,
    48'h0000000df8640,
    48'h0000000df8641,
    48'h0000000df8642,
    48'h0000000df8643,
    48'h0000000df8644,
    48'h0000000df8645,
    48'h0000000df8646,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df8648,
    48'h0000000df8649,
    48'h0000040138938,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034d71,
    48'h0000040138938,
    48'h0000040138940,
    48'h0000042354e20,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h000007b034d72,
    48'h0000000df864a,
    48'h0000000df864b,
    48'h0000040138938,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034d71,
    48'h0000040138938,
    48'h0000040138940,
    48'h0000042354e20,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h000007b034d72,
    48'h0000000df864c,
    48'h0000000df864d,
    48'h0000000df864e,
    48'h0000000df864f,
    48'h0000000df8650,
    48'h0000000df8651,
    48'h0000000df8652,
    48'h0000040138940,
    48'h000007b034d98,
    48'h000007b034c70,
    48'h0000000df8654,
    48'h0000000df8655,
    48'h0000000df8656,
    48'h0000000df8657,
    48'h0000000df8658,
    48'h0000000df8659,
    48'h0000000df865a,
    48'h0000000df865b,
    48'h0000000df865c,
    48'h0000000df865d,
    48'h0000000df865e,
    48'h0000000df865f,
    48'h0000000df8660,
    48'h0000000df8661,
    48'h0000000df8662,
    48'h0000000df8663,
    48'h0000000df8664,
    48'h0000000df8665,
    48'h0000000df8666,
    48'h0000040138938,
    48'h0000042354e20,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df863c,
    48'h0000040138938,
    48'h0000042354e24,
    48'h00000401367d0,
    48'h000007b0345b4,
    48'h0000040136428,
    48'h000007b034a34,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df8648,
    48'h000004013893c,
    48'h0000042354e24,
    48'h00000401367d0,
    48'h000007b0345b4,
    48'h0000040136428,
    48'h000007b034a34,
    48'h0000040138940,
    48'h0000042351e00,
    48'h000007b034d60,
    48'h000007b034c88,
    48'h000007b034c70,
    48'h0000000df8654,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354e20,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df863c,
    48'h0000000df863c,
    48'h000007b034d58,
    48'h0000000df863d,
    48'h000007b034dfc,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000000df863e,
    48'h000007b034c68,
    48'h000007b034cc0,
    48'h000007b034cb8,
    48'h000007b034de4,
    48'h0000042354e20,
    48'h000007b034c98,
    48'h000007b034cc8,
    48'h000007b034de4,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df8648,
    48'h0000000df8648,
    48'h0000000df8649,
    48'h000007b034ccc,
    48'h000007b034ddc,
    48'h000007b034d71,
    48'h000007b034cb0,
    48'h000007b034c98,
    48'h000007b034c9c,
    48'h0000000df864a,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034cb9,
    48'h0000042354e20,
    48'h000007b034c9c,
    48'h000007b034ccc,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h0000042351e00,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df8654,
    48'h0000000df8654,
    48'h000007b034ca0,
    48'h0000040139a84,
    48'h000007b034ca0,
    48'h0000042351e00,
    48'h0000000df8655,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df8656,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df8657,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df8658,
    48'h0000042351e00,
    48'h0000000df8659,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034dfc,
    48'h000007b034cb2,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034dec,
    48'h000007b034de4,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354e20,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df863f,
    48'h0000000df863f,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354e20,
    48'h0000040138938,
    48'h0000042354e22,
    48'h000007b034c98,
    48'h0000042354e24,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df8640,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df864b,
    48'h0000000df864b,
    48'h000007b034ccc,
    48'h000007b034ddc,
    48'h000007b034d71,
    48'h000007b034cb0,
    48'h000007b034c98,
    48'h000007b034c9c,
    48'h0000000df864c,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h0000042351e00,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df865a,
    48'h0000000df865a,
    48'h000007b034dfc,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000000df865b,
    48'h000007b034ca0,
    48'h0000040139a98,
    48'h000007b034ca0,
    48'h0000042351e00,
    48'h0000000df865c,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df865d,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df865e,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df865f,
    48'h0000042351e00,
    48'h0000000df8660,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034dfc,
    48'h000007b034cb2,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034d94,
    48'h000004013893c,
    48'h000007b034d98,
    48'h0000040138940,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034d42,
    48'h000007b034ca0,
    48'h000007b034ce8,
    48'h000007b034cba,
    48'h000007b034d4a,
    48'h000007b034cd0,
    48'h000007b034d18,
    48'h000007b034cc2,
    48'h000007b034d52,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d30,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d42,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423afd84,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423afd74,
    48'h000007b034cfc,
    48'h0000040139dd8,
    48'h000007b034d98,
    48'h00000423afd78,
    48'h000007b034d00,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d42,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e20,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h000007b034d42,
    48'h000007b034d30,
    48'h000007b034d18,
    48'h00000400015a4,
    48'h0000040138940,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8124,
    48'h0000040136800,
    48'h00000423afdb4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423ae428,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423ae438,
    48'h00000423ae418,
    48'h00000423ae41c,
    48'h0000042351df0,
    48'h00000423ae418,
    48'h00000423ae418,
    48'h00000423ae420,
    48'h0000042354d90,
    48'h00000423ae418,
    48'h000004214c8a8,
    48'h00000423ae43c,
    48'h00000423ae43c,
    48'h000007b034dcc,
    48'h0000000dfcf34,
    48'h000007b034dd4,
    48'h0000000df7bd4,
    48'h000007b034dd4,
    48'h00000423ae43c,
    48'h00000423ae438,
    48'h00000423ae43c,
    48'h00000400025c0,
    48'h0000040139dd0,
    48'h00000423ae420,
    48'h0000040138938,
    48'h000007b034dcc,
    48'h0000000df882c,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9ccc,
    48'h000007b034da8,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df8420,
    48'h0000000df8421,
    48'h0000000df8422,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df8420,
    48'h0000040138938,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040136428,
    48'h000007b034a50,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df8420,
    48'h0000000df8420,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354d90,
    48'h0000040138938,
    48'h0000042354d92,
    48'h000007b034c98,
    48'h0000042354d94,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df8421,
    48'h000007b034dfc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000000df8422,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034cc0,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d40,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423ae420,
    48'h000007b034cf8,
    48'h000007b034d40,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d90,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df7ff4,
    48'h0000040136800,
    48'h00000423ae434,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423ae498,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423ae4a8,
    48'h00000423ae488,
    48'h00000423ae48c,
    48'h0000042351de8,
    48'h00000423ae488,
    48'h00000423ae488,
    48'h00000423ae490,
    48'h00000423ae478,
    48'h00000423ae488,
    48'h000004214c8a8,
    48'h00000423ae4ac,
    48'h00000423ae4ac,
    48'h000007b034dcc,
    48'h0000000dfd28c,
    48'h000007b034dd4,
    48'h0000000df7f2c,
    48'h000007b034dd4,
    48'h0000040136800,
    48'h00000423ae4a4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423afe90,
    48'h00000423afe90,
    48'h00000423afe9c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423b0050,
    48'h00000423b0050,
    48'h00000423b005c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2d0,
    48'h00000423afeb8,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afec8,
    48'h00000423afea8,
    48'h00000423afeac,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h00000423afeb0,
    48'h0000042351e00,
    48'h00000423afea8,
    48'h00000423afea8,
    48'h00000423afeb0,
    48'h0000042351e00,
    48'h00000423afea8,
    48'h000004214c8a8,
    48'h00000423afecc,
    48'h00000423afecc,
    48'h000007b034dcc,
    48'h0000000dfcfa8,
    48'h000007b034dd4,
    48'h0000000df7c48,
    48'h000007b034dd4,
    48'h00000423afecc,
    48'h00000423afec8,
    48'h00000423afecc,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423afeac,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423afeb0,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df8a70,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9f10,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8a74,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000df9f14,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354c70,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354c74,
    48'h00000401367d0,
    48'h000007b0345a8,
    48'h0000040136428,
    48'h000007b034a28,
    48'h000004013893c,
    48'h0000042351e00,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354c70,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b034d58,
    48'h0000000df84d5,
    48'h000007b034dfc,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354c70,
    48'h0000040138938,
    48'h0000042354c72,
    48'h000007b034c98,
    48'h0000042354c74,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e00,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034c9c,
    48'h0000040139a84,
    48'h000007b034c9c,
    48'h0000042351e00,
    48'h0000000df84e5,
    48'h000007b034c9c,
    48'h0000040139bac,
    48'h000007b034c9c,
    48'h0000042351e00,
    48'h0000000df84e6,
    48'h000007b034c9c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034c9c,
    48'h0000042351e00,
    48'h0000000df84e7,
    48'h000007b034dfc,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000000df84e8,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df84e9,
    48'h0000042351e00,
    48'h0000000df84ea,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034cb9,
    48'h0000042351e00,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034dec,
    48'h000007b034de4,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb0,
    48'h000007b034d40,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb1,
    48'h000007b034d41,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354c70,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d7,
    48'h0000000df84d7,
    48'h000007b034c98,
    48'h0000040139a84,
    48'h000007b034c98,
    48'h0000042354c70,
    48'h0000040138938,
    48'h0000042354c72,
    48'h000007b034c98,
    48'h0000042354c74,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df84d8,
    48'h000007b034c98,
    48'h0000040139bac,
    48'h000007b034c98,
    48'h0000042354c70,
    48'h0000040138938,
    48'h0000042354c72,
    48'h000007b034c98,
    48'h0000042354c74,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d9,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e00,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84eb,
    48'h0000000df84eb,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000000df84ec,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423afeac,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423afeb0,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h0000042354c70,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8068,
    48'h0000040136800,
    48'h00000423afec4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2d0,
    48'h00000423afee0,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afef0,
    48'h00000423afed8,
    48'h0000040136800,
    48'h00000423afeec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2d0,
    48'h00000423aff58,
    48'h00000423aff58,
    48'h00000423aff64,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2d0,
    48'h0000042354c78,
    48'h0000042354c78,
    48'h0000042354c84,
    48'h000007b0343c8,
    48'h000007b0343cc,
    48'h000007b0343d0,
    48'h000007b0343d4,
    48'h000007b0343d8,
    48'h000007b0343dc,
    48'h000007b0343e0,
    48'h000007b0343e4,
    48'h000007b0343e8,
    48'h000007b0343ec,
    48'h000007b0343f0,
    48'h000007b0343f4,
    48'h000007b0343f8,
    48'h000007b0343fc,
    48'h0000040023890,
    48'h000007b034390,
    48'h000007b034400,
    48'h000007b034438,
    48'h000007b034394,
    48'h000007b034404,
    48'h000007b03443c,
    48'h000007b034398,
    48'h000007b034408,
    48'h000007b034440,
    48'h000007b03439c,
    48'h000007b03440c,
    48'h000007b034444,
    48'h000007b0343a0,
    48'h000007b034410,
    48'h000007b034448,
    48'h000007b0343a4,
    48'h000007b034524,
    48'h0000040023890,
    48'h000007b034400,
    48'h000007b034390,
    48'h000007b034438,
    48'h000007b034404,
    48'h000007b034394,
    48'h000007b03443c,
    48'h000007b034408,
    48'h000007b034398,
    48'h000007b034440,
    48'h000007b03440c,
    48'h000007b03439c,
    48'h000007b034444,
    48'h000007b034410,
    48'h000007b0343a0,
    48'h000007b034448,
    48'h000007b034414,
    48'h000007b0343a4,
    48'h0000040023b70,
    48'h0000040002490,
    48'h000007b034c14,
    48'h000007b034c10,
    48'h0000040023b70,
    48'h000007b034c10,
    48'h0000040023b70,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040023892,
    48'h0000040023a5a,
    48'h0000040023aca,
    48'h000007b0343a4,
    48'h000007b0343a4,
    48'h0000040139780,
    48'h0000040139780,
    48'h000007b0343a8,
    48'h000007b0343a8,
    48'h0000040139784,
    48'h0000040139784,
    48'h000007b0343ac,
    48'h000007b0343ac,
    48'h0000040139788,
    48'h0000040139788,
    48'h000007b0343b0,
    48'h000007b0343b0,
    48'h000004013978c,
    48'h000004013978c,
    48'h000007b0343b8,
    48'h000007b0343b8,
    48'h0000040139790,
    48'h0000040139790,
    48'h000007b0343bc,
    48'h000007b0343bc,
    48'h0000040139794,
    48'h0000040139794,
    48'h000007b0343c0,
    48'h000007b0343c0,
    48'h0000040139798,
    48'h0000040139798,
    48'h000007b0343c4,
    48'h000007b0343c4,
    48'h000004013979c,
    48'h000007b03444c,
    48'h000007b034c14,
    48'h0000040023890,
    48'h0000040023b38,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc0,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc2,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc4,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc6,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc8,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbca,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbcc,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbce,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd0,
    48'h0000040139068,
    48'h0000042352bd0,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd2,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd4,
    48'h0000040139068,
    48'h0000042352bd8,
    48'h00000423ace3a,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd6,
    48'h0000040139068,
    48'h0000042352bdc,
    48'h00000423aceca,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd8,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbda,
    48'h0000040139068,
    48'h0000042352be4,
    48'h00000423ad2ca,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbdc,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbde,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe0,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe2,
    48'h0000040139068,
    48'h0000042352bf4,
    48'h00000423adaea,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe4,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe6,
    48'h0000040139068,
    48'h0000042352bfc,
    48'h00000423ae05a,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe8,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbea,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbec,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbee,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbf0,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbf2,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbf4,
    48'h000004214c578,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040023890,
    48'h0000040138b29,
    48'h000007b0343a4,
    48'h000007b03444c,
    48'h000007b034418,
    48'h000007b0343a8,
    48'h000007b034450,
    48'h000007b03441c,
    48'h000007b0343ac,
    48'h000007b034454,
    48'h000007b034420,
    48'h000007b0343b0,
    48'h000007b034458,
    48'h000007b034424,
    48'h000007b0343b4,
    48'h000007b03445c,
    48'h000007b034428,
    48'h000007b0343b8,
    48'h000007b034460,
    48'h000007b03442c,
    48'h000007b0343bc,
    48'h000007b034464,
    48'h000007b034430,
    48'h000007b0343c0,
    48'h000007b034468,
    48'h000007b034434,
    48'h000007b0343c4,
    48'h000007b03446c,
    48'h000004213c268,
    48'h0000040139038,
    48'h000007b03451c,
    48'h000004214c578,
    48'h0000040023760,
    48'h000004214c578,
    48'h0000040023768,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h0000042354b84,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354b78,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354b7a,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h0000042354b88,
    48'h0000042354b68,
    48'h0000042354b6c,
    48'h0000042354b60,
    48'h0000042354b64,
    48'h0000042354b70,
    48'h0000042354af8,
    48'h0000042354b68,
    48'h0000042354b68,
    48'h0000042354b70,
    48'h0000042354af8,
    48'h0000042354b68,
    48'h000004214c8a8,
    48'h0000042354b8c,
    48'h0000042354b8c,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h0000042354b8c,
    48'h0000042354b88,
    48'h0000042354b8c,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h0000042354b6c,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042354b70,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354b60,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354b64,
    48'h00000401367d0,
    48'h000007b0345c0,
    48'h0000040136428,
    48'h000007b034a40,
    48'h000004013893c,
    48'h0000042354af8,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h0000042354afa,
    48'h0000042354afc,
    48'h0000042354ae8,
    48'h0000042354ae8,
    48'h0000042354ae8,
    48'h0000042354ae8,
    48'h0000042354ae8,
    48'h0000042354aec,
    48'h0000042351e40,
    48'h0000042351e44,
    48'h0000042354af0,
    48'h0000042354ae0,
    48'h0000042354ae4,
    48'h0000042354ae8,
    48'h0000042354af0,
    48'h0000042354ae0,
    48'h0000042354aec,
    48'h0000042351e40,
    48'h0000042351e44,
    48'h00000401367d0,
    48'h000007b0345e0,
    48'h0000040139dd4,
    48'h0000042354b70,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042354b60,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042354b60,
    48'h0000042354b64,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042354b60,
    48'h0000040138938,
    48'h0000042354b62,
    48'h000007b034f58,
    48'h0000042354b64,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042354af8,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042354af8,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042354af8,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042354af8,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000000df84e8,
    48'h0000042354af8,
    48'h0000000df84e9,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h0000042354b6c,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042354b70,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354b60,
    48'h0000042354b60,
    48'h0000042354b64,
    48'h0000042354b60,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354afa,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042354b70,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042354b70,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034ba8,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000042354b88,
    48'h0000042354b68,
    48'h0000042354b6c,
    48'h0000042354b60,
    48'h0000042354b60,
    48'h0000042354b60,
    48'h0000042354b64,
    48'h0000042354b62,
    48'h0000040001fac,
    48'h0000040023a64,
    48'h0000040023768,
    48'h000007b034e2e,
    48'h0000040023760,
    48'h000007b034cc0,
    48'h0000042354b94,
    48'h0000042354b9a,
    48'h0000042354ba0,
    48'h0000042354b78,
    48'h0000042354b78,
    48'h000004213c310,
    48'h0000042354c4c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354c40,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354c42,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h0000042354c50,
    48'h0000042354c30,
    48'h0000042354c34,
    48'h0000042354c28,
    48'h0000042354c2c,
    48'h0000042354c38,
    48'h0000042354bc0,
    48'h0000042354c30,
    48'h0000042354c30,
    48'h0000042354c38,
    48'h0000042354bc0,
    48'h0000042354c30,
    48'h000004214c8a8,
    48'h0000042354c54,
    48'h0000042354c54,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h0000042354c54,
    48'h0000042354c50,
    48'h0000042354c54,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h0000042354c34,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042354c38,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354c28,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354c2c,
    48'h00000401367d0,
    48'h000007b0345bc,
    48'h0000040136428,
    48'h000007b034a3c,
    48'h000004013893c,
    48'h0000042354bc0,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h0000042354bc2,
    48'h0000042354bc4,
    48'h0000042354bb0,
    48'h0000042354bb0,
    48'h0000042354bb0,
    48'h0000042354bb0,
    48'h0000042354bb0,
    48'h0000042354bb4,
    48'h0000042351e40,
    48'h0000042351e44,
    48'h0000042354bb8,
    48'h0000042354ba8,
    48'h0000042354bac,
    48'h0000042354bb0,
    48'h0000042354bb8,
    48'h0000042354ba8,
    48'h0000042354bb4,
    48'h0000042351e40,
    48'h0000042351e44,
    48'h00000401367d0,
    48'h000007b0345e0,
    48'h0000040139dd4,
    48'h0000042354c38,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042354c28,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042354c28,
    48'h0000042354c2c,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042354c28,
    48'h0000040138938,
    48'h0000042354c2a,
    48'h000007b034f58,
    48'h0000042354c2c,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042354bc0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042354bc0,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042354bc0,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042354bc0,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000000df84e8,
    48'h0000042354bc0,
    48'h0000000df84e9,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h0000042354c34,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042354c38,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354c28,
    48'h0000042354c28,
    48'h0000042354c2c,
    48'h0000042354c28,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042354c38,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042354c38,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034ba8,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000042354c50,
    48'h0000042354c30,
    48'h0000042354c34,
    48'h0000042354c28,
    48'h0000042354c28,
    48'h0000042354c28,
    48'h0000042354c2c,
    48'h0000042354c2a,
    48'h0000040001fac,
    48'h0000040023a62,
    48'h0000040023768,
    48'h000007b034e2d,
    48'h0000040023760,
    48'h000007b034cbc,
    48'h0000042354c5c,
    48'h0000042354c62,
    48'h0000042354c68,
    48'h0000042354c40,
    48'h0000042354c40,
    48'h000004213c310,
    48'h0000042354c9c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354c90,
    48'h0000042354c90,
    48'h0000042354c90,
    48'h0000042354c90,
    48'h000004213c310,
    48'h0000042354d24,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354d18,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354d1a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042354d28,
    48'h0000042354d08,
    48'h0000042354d0c,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042354d02,
    48'h0000040001fac,
    48'h0000040023a6e,
    48'h0000040023768,
    48'h000007b034e33,
    48'h0000040023760,
    48'h000007b034cd4,
    48'h0000042354d34,
    48'h0000042354d18,
    48'h0000042354d18,
    48'h000004213c310,
    48'h0000042354db4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354da8,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354daa,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042354db8,
    48'h0000042354d98,
    48'h0000042354d9c,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d92,
    48'h0000040001fac,
    48'h0000040023a6c,
    48'h0000040023768,
    48'h000007b034e32,
    48'h0000040023760,
    48'h000007b034cd0,
    48'h0000042354dc4,
    48'h0000042354da8,
    48'h0000042354da8,
    48'h000004213c310,
    48'h0000042354ebc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354eb0,
    48'h0000042354eb0,
    48'h0000042354eb0,
    48'h0000042354eb0,
    48'h000004213c310,
    48'h0000042354eec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354ee0,
    48'h0000042354ee0,
    48'h0000042354ee0,
    48'h0000042354ee0,
    48'h000004213c310,
    48'h0000042354f1c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354f10,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354f12,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042354f20,
    48'h0000042354f00,
    48'h0000042354f04,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h0000040023a5e,
    48'h0000040023768,
    48'h000007b034e2b,
    48'h0000040023760,
    48'h000007b034cb4,
    48'h0000042354f2c,
    48'h0000042354f10,
    48'h0000042354f10,
    48'h000004213c310,
    48'h00000423b032c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h00000423b0320,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423b0322,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423b0330,
    48'h00000423b0310,
    48'h00000423b0314,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h00000423b033c,
    48'h00000423b0320,
    48'h00000423b0320,
    48'h000004213c310,
    48'h00000423b03a4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h00000423b0398,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423b039a,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423b03a8,
    48'h00000423b0358,
    48'h00000423b035c,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h00000423b03b4,
    48'h00000423b0398,
    48'h00000423b0398,
    48'h000004213c310,
    48'h0000042354f6c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354f60,
    48'h0000042354f60,
    48'h0000042354f60,
    48'h0000042354f60,
    48'h000004213c310,
    48'h00000423557a4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042355798,
    48'h0000042355798,
    48'h0000042355798,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042355798,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h0000042355054,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af260,
    48'h0000042355048,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235504a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042355064,
    48'h0000042355048,
    48'h0000042355048,
    48'h000004213c310,
    48'h00000423550c4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af260,
    48'h00000423550b8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423550ba,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423550c8,
    48'h00000423550a8,
    48'h00000423550ac,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h00000423550d4,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h000004213c310,
    48'h00000423550ec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af260,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h000004213c310,
    48'h000004235515c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af260,
    48'h0000042355150,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355152,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h000004235513c,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355140,
    48'h0000042355140,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355140,
    48'h000004214c8a8,
    48'h0000042355164,
    48'h0000042355164,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h0000042355164,
    48'h0000042355160,
    48'h0000042355164,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h0000042355144,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042355148,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042355138,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h000004235513c,
    48'h00000401367d0,
    48'h000007b0345c8,
    48'h0000040136428,
    48'h000007b034a48,
    48'h000004013893c,
    48'h0000042355130,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h0000042355132,
    48'h0000042355134,
    48'h0000042355120,
    48'h0000042355120,
    48'h0000042355120,
    48'h0000042355120,
    48'h0000042355120,
    48'h0000042355124,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042355128,
    48'h0000042355118,
    48'h000004235511c,
    48'h0000042355120,
    48'h0000042355128,
    48'h0000042355118,
    48'h0000042355124,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040139dd4,
    48'h0000042355148,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355138,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042355138,
    48'h000004235513c,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042355138,
    48'h0000040138938,
    48'h000004235513a,
    48'h000007b034f58,
    48'h000004235513c,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042355130,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042355130,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042355130,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042355130,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000000df84e8,
    48'h0000042355130,
    48'h0000000df84e9,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h0000042355144,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042355148,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042355138,
    48'h0000042355138,
    48'h000004235513c,
    48'h0000042355138,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355130,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355132,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042355148,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042355148,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034baa,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c780,
    48'h0000040139978,
    48'h000004214c490,
    48'h0000042355130,
    48'h0000040138f40,
    48'h0000042355130,
    48'h000004214c490,
    48'h0000040139978,
    48'h000004214c698,
    48'h0000042355130,
    48'h0000042355130,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c490,
    48'h0000040139540,
    48'h000007b035194,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355134,
    48'h0000042355130,
    48'h0000042355120,
    48'h00000400015bc,
    48'h0000042355158,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e8,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h00000423550c0,
    48'h0000042355048,
    48'h0000042355048,
    48'h000007b035154,
    48'h000004235504c,
    48'h000004213a120,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042355040,
    48'h0000042354d90,
    48'h000004235503c,
    48'h0000042355130,
    48'h0000042351df0,
    48'h0000042355050,
    48'h0000042355798,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000007b034fb8,
    48'h0000040139978,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h0000042355138,
    48'h0000042355138,
    48'h000004235513c,
    48'h000004235513a,
    48'h0000040001fac,
    48'h0000040023a68,
    48'h0000040023768,
    48'h000007b034e30,
    48'h0000040023760,
    48'h000007b034cc8,
    48'h000004235516c,
    48'h0000042355150,
    48'h0000042355150,
    48'h000004213c310,
    48'h00000423551ec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af264,
    48'h00000423551e0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423551e2,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423551f0,
    48'h00000423551d0,
    48'h00000423551d4,
    48'h0000042351df0,
    48'h00000423551d0,
    48'h00000423551d0,
    48'h00000423551d8,
    48'h00000423551c0,
    48'h00000423551d0,
    48'h000004214c8a8,
    48'h00000423551f4,
    48'h00000423551f4,
    48'h000007b03508c,
    48'h0000000dfcf58,
    48'h000007b035094,
    48'h0000000df7bf8,
    48'h000007b035094,
    48'h00000423551f4,
    48'h00000423551f0,
    48'h00000423551f4,
    48'h00000400025e4,
    48'h00000423551d8,
    48'h0000040139dd0,
    48'h00000423551c4,
    48'h0000040138938,
    48'h00000423551d8,
    48'h0000040139dd4,
    48'h00000423551c8,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df88e0,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9d80,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df88e4,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9d84,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df8444,
    48'h0000000df8445,
    48'h0000000df8446,
    48'h0000000df8447,
    48'h0000000df8448,
    48'h0000000df8449,
    48'h0000000df844a,
    48'h0000000df844b,
    48'h0000000df844c,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df8450,
    48'h0000000df8451,
    48'h0000000df8452,
    48'h0000000df8453,
    48'h0000000df8454,
    48'h0000000df8455,
    48'h0000000df8456,
    48'h0000000df8457,
    48'h0000000df8458,
    48'h0000040138938,
    48'h0000042355190,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df8444,
    48'h0000040138938,
    48'h0000040139dd0,
    48'h0000042355192,
    48'h0000042355194,
    48'h0000042355180,
    48'h0000042355180,
    48'h0000042355180,
    48'h0000042355180,
    48'h0000042355180,
    48'h0000042355184,
    48'h0000042355138,
    48'h000004235513c,
    48'h0000042355188,
    48'h0000042355178,
    48'h000004235517c,
    48'h0000042355180,
    48'h0000042355188,
    48'h0000042355178,
    48'h0000042355184,
    48'h0000042355138,
    48'h000004235513c,
    48'h00000401367d0,
    48'h000007b0345c8,
    48'h0000040139dd0,
    48'h00000423551c4,
    48'h0000040138938,
    48'h000007b035050,
    48'h000004013893c,
    48'h00000423551b8,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df8450,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423551ba,
    48'h00000423551bc,
    48'h00000423551a8,
    48'h00000423551a8,
    48'h00000423551a8,
    48'h00000423551a8,
    48'h00000423551a8,
    48'h00000423551ac,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423551b0,
    48'h00000423551a0,
    48'h00000423551a4,
    48'h00000423551a8,
    48'h00000423551b0,
    48'h00000423551a0,
    48'h00000423551ac,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h00000423551c8,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355190,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df8444,
    48'h0000000df8444,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042355190,
    48'h0000000df8445,
    48'h0000042355190,
    48'h0000000df8446,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000000df8447,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h0000042355190,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423551b8,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8450,
    48'h0000000df8450,
    48'h000007b0350bc,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h0000000df8451,
    48'h000007b034f5c,
    48'h0000040139a98,
    48'h000007b034f5c,
    48'h00000423551b8,
    48'h0000000df8452,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355190,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df8448,
    48'h0000000df8448,
    48'h000007b0350bc,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000000df8449,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042355190,
    48'h0000000df844a,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423551b8,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8453,
    48'h0000000df8453,
    48'h00000423551b8,
    48'h0000000df8454,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h0000000df8455,
    48'h000007b034f5c,
    48'h0000040139a98,
    48'h000007b034f5c,
    48'h00000423551b8,
    48'h0000000df8456,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423551b8,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355190,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df844b,
    48'h0000000df844b,
    48'h0000042355190,
    48'h000007b034f40,
    48'h0000042355194,
    48'h0000042355180,
    48'h0000000df844c,
    48'h000007b034f28,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h000007b0350a4,
    48'h0000042355190,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423551b8,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8457,
    48'h0000000df8457,
    48'h00000423551b8,
    48'h000007b034f44,
    48'h00000423551bc,
    48'h00000423551a8,
    48'h0000000df8458,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h000007b0350a4,
    48'h00000423551b8,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b034fd0,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423551c4,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423551c8,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h0000040138938,
    48'h0000042355190,
    48'h0000042355190,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fd0,
    48'h000007b034fe8,
    48'h000007b035008,
    48'h000007b034fe8,
    48'h000007b035018,
    48'h0000040138938,
    48'h000007b035018,
    48'h000007b034fa0,
    48'h000007b035154,
    48'h000007b035018,
    48'h000007b035068,
    48'h000007b035150,
    48'h000007b035018,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb17b,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd0,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355192,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423551c4,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423551c4,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fb8,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb17c,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551ba,
    48'h0000040136800,
    48'h0000040139540,
    48'h000004214c780,
    48'h000004214c490,
    48'h0000042355190,
    48'h0000042355190,
    48'h00000423551b8,
    48'h0000042355192,
    48'h00000423551ba,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h0000042355194,
    48'h00000423551bc,
    48'h0000042355180,
    48'h00000423551a8,
    48'h0000042355182,
    48'h00000423551aa,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h0000042355188,
    48'h00000423551b0,
    48'h0000042355178,
    48'h00000423551a0,
    48'h000004235517a,
    48'h00000423551a2,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h000004235517c,
    48'h00000423551a4,
    48'h00000003840fc,
    48'h0000042355184,
    48'h00000423551ac,
    48'h0000042355138,
    48'h0000042354d90,
    48'h000004235513a,
    48'h0000042354d92,
    48'h000004235513c,
    48'h0000042354d94,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040139540,
    48'h000004214c780,
    48'h000004214c698,
    48'h00000423551b8,
    48'h000004214c490,
    48'h0000042355190,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c494,
    48'h000004214c69c,
    48'h0000040139544,
    48'h000004214c344,
    48'h000004013885c,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136514,
    48'h000004214c781,
    48'h000004214c599,
    48'h00000423551c8,
    48'h0000040136800,
    48'h0000040138f44,
    48'h00000423551c8,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h0000040022cc4,
    48'h0000040022de8,
    48'h0000040022ccc,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000004214c69c,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8018,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034baa,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000007b034ff4,
    48'h000004214c344,
    48'h000004013885c,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c344,
    48'h0000040139544,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h0000040021af0,
    48'h0000040021af8,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h0000040138eb0,
    48'h0000040138eb1,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h0000040138eb0,
    48'h0000040138eb1,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c780,
    48'h0000040139978,
    48'h000004214c490,
    48'h0000042355190,
    48'h0000040138f40,
    48'h0000042355190,
    48'h000004214c490,
    48'h0000040139978,
    48'h000004214c698,
    48'h0000042355190,
    48'h0000042355190,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c490,
    48'h0000040139540,
    48'h000007b035194,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355194,
    48'h0000042355190,
    48'h0000042355180,
    48'h00000400015bc,
    48'h00000423551e8,
    48'h0000042355150,
    48'h0000042355150,
    48'h000007b035154,
    48'h0000042355154,
    48'h000004213a120,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h0000042355148,
    48'h0000042355190,
    48'h0000042355130,
    48'h0000042355192,
    48'h0000042355132,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h0000042355194,
    48'h0000042355134,
    48'h0000042355180,
    48'h0000042355120,
    48'h0000042355182,
    48'h0000042355122,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h0000042355188,
    48'h0000042355128,
    48'h0000042355178,
    48'h0000042355118,
    48'h000004235517c,
    48'h000004235511c,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355158,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e8,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h00000423550c0,
    48'h0000042355048,
    48'h0000042355048,
    48'h000007b035154,
    48'h000004235504c,
    48'h000004213a120,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042355040,
    48'h0000042354d90,
    48'h000004235503c,
    48'h0000042355190,
    48'h0000042351df0,
    48'h0000042355050,
    48'h0000042355798,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040023890,
    48'h0000040023b38,
    48'h000007b034f11,
    48'h0000040139540,
    48'h0000040023b38,
    48'h00000400024b8,
    48'h0000040023b38,
    48'h0000040001fac,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040001fac,
    48'h0000040023b38,
    48'h000007b034f11,
    48'h0000040023b38,
    48'h0000040023a5a,
    48'h00000400237b0,
    48'h0000040023898,
    48'h0000040023b38,
    48'h000007b035158,
    48'h000007b03515c,
    48'h000007b035160,
    48'h000007b035164,
    48'h000007b035164,
    48'h000007b035160,
    48'h000004214c960,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b09e0,
    48'h00000423b09e0,
    48'h00000423b09e2,
    48'h0000040002104,
    48'h000004214c960,
    48'h0000000384108,
    48'h000007b03515c,
    48'h00000423b09e4,
    48'h000004214c960,
    48'h0000040023898,
    48'h0000040139978,
    48'h000007b034ff0,
    48'h0000040139978,
    48'h00000423b09e4,
    48'h00000401364c8,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000004214c344,
    48'h000004214c69c,
    48'h000004214c494,
    48'h000004013885c,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c781,
    48'h000004013997c,
    48'h000004214c494,
    48'h00000423551b8,
    48'h0000040138f44,
    48'h00000423551b8,
    48'h000004214c494,
    48'h000004013997c,
    48'h000004214c69c,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c494,
    48'h0000040139544,
    48'h000007b035194,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551bc,
    48'h00000423551b8,
    48'h00000423551a8,
    48'h00000400015bc,
    48'h00000423551e8,
    48'h0000042355150,
    48'h0000042355150,
    48'h000007b035154,
    48'h0000042355154,
    48'h000004213a120,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h0000042355148,
    48'h00000423551b8,
    48'h0000042355130,
    48'h00000423551ba,
    48'h0000042355132,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h00000423551bc,
    48'h0000042355134,
    48'h00000423551a8,
    48'h0000042355120,
    48'h00000423551aa,
    48'h0000042355122,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h00000423551b0,
    48'h0000042355128,
    48'h00000423551a0,
    48'h0000042355118,
    48'h00000423551a4,
    48'h000004235511c,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355158,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e8,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h00000423550c0,
    48'h0000042355048,
    48'h0000042355048,
    48'h000007b035154,
    48'h000004235504c,
    48'h000004213a120,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042355040,
    48'h0000042354d90,
    48'h000004235503c,
    48'h00000423551b8,
    48'h0000042351df0,
    48'h0000042355050,
    48'h0000042355798,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h0000040139978,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000042355190,
    48'h0000040138f40,
    48'h0000042355190,
    48'h00000400237b0,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000007b034ff4,
    48'h000004214c69c,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000007b034fb8,
    48'h0000040139978,
    48'h0000042355192,
    48'h000004214c780,
    48'h0000042355190,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035194,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355194,
    48'h0000042355190,
    48'h0000042355180,
    48'h00000400015bc,
    48'h00000423551e8,
    48'h0000042355150,
    48'h0000042355150,
    48'h000007b035154,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h0000042355148,
    48'h0000042355190,
    48'h0000042355130,
    48'h0000042355192,
    48'h0000042355132,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h0000042355194,
    48'h0000042355134,
    48'h0000042355180,
    48'h0000042355120,
    48'h0000042355182,
    48'h0000042355122,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h0000042355188,
    48'h0000042355128,
    48'h0000042355178,
    48'h0000042355118,
    48'h000004235517c,
    48'h000004235511c,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355158,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e8,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h00000423550c0,
    48'h0000042355048,
    48'h0000042355048,
    48'h000007b035154,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042355040,
    48'h0000042354d90,
    48'h000004235503c,
    48'h0000042355190,
    48'h0000042351df0,
    48'h0000042355050,
    48'h0000042355798,
    48'h00000423b09e2,
    48'h0000042355190,
    48'h0000042355192,
    48'h0000042355190,
    48'h00000400015a4,
    48'h0000042355190,
    48'h00000423b09e2,
    48'h000004213a240,
    48'h000004235914c,
    48'h0000000df7828,
    48'h000007b035258,
    48'h000007b03525c,
    48'h000007b035260,
    48'h000007b035264,
    48'h000007b035264,
    48'h000007b035260,
    48'h000004214c93c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b09e8,
    48'h00000423b09e8,
    48'h00000423b09ea,
    48'h00000400020e0,
    48'h000004214c93c,
    48'h00000003840fc,
    48'h000007b03525c,
    48'h00000423b09ec,
    48'h000004214c93c,
    48'h00000003840fd,
    48'h000007b035258,
    48'h00000423b09f0,
    48'h000004214c93c,
    48'h00000423b09e8,
    48'h000004214c90c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b09f8,
    48'h00000423b09f8,
    48'h00000423b0a0c,
    48'h00000423b0a10,
    48'h00000423b0a08,
    48'h00000423b0a14,
    48'h0000040002394,
    48'h0000040002394,
    48'h00000423b09fc,
    48'h00000423551e8,
    48'h00000423b0a04,
    48'h00000423b0a00,
    48'h00000423b0a00,
    48'h000004235515c,
    48'h00000423551e8,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040023978,
    48'h0000040136800,
    48'h000004214c494,
    48'h000007b034fb9,
    48'h000004013997c,
    48'h00000400015a4,
    48'h000007b034fb9,
    48'h000004214c69c,
    48'h000007b034ff4,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h00000423b09e2,
    48'h0000040022cc0,
    48'h0000040022cb8,
    48'h00000423551c4,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h000004013997c,
    48'h0000040022cc8,
    48'h0000040138eb1,
    48'h0000040022de8,
    48'h00000423551f0,
    48'h00000423551d0,
    48'h00000423551d4,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h00000423551fc,
    48'h00000423b03f2,
    48'h00000423b03f8,
    48'h00000423551e0,
    48'h00000423551e0,
    48'h000004213c310,
    48'h000004235525c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af264,
    48'h0000042355250,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355252,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355260,
    48'h0000042355240,
    48'h0000042355244,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235526c,
    48'h0000042355250,
    48'h0000042355250,
    48'h000004213c310,
    48'h0000042355294,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af264,
    48'h0000042355288,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235528a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355298,
    48'h0000042355278,
    48'h000004235527c,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h0000042354c72,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h0000040023760,
    48'h000007b034ca8,
    48'h00000423552a4,
    48'h0000042355288,
    48'h0000042355288,
    48'h000004213c310,
    48'h00000423552bc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af268,
    48'h00000423552b0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423552b2,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423552c0,
    48'h00000423552a8,
    48'h00000423552a8,
    48'h00000423552cc,
    48'h00000423b0412,
    48'h00000423b0418,
    48'h00000423552b0,
    48'h00000423552b0,
    48'h000004213c310,
    48'h00000423552fc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af268,
    48'h00000423552f0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423552f2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355300,
    48'h00000423552e0,
    48'h00000423552e4,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235530c,
    48'h00000423552f0,
    48'h00000423552f0,
    48'h000004213c310,
    48'h0000042355324,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af268,
    48'h0000042355318,
    48'h0000042355318,
    48'h0000042355318,
    48'h0000042355318,
    48'h000004213c310,
    48'h0000042355104,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af268,
    48'h00000423550f8,
    48'h00000423550f8,
    48'h00000423550f8,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h00000423550f8,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423553a4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af26c,
    48'h0000042355398,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235539a,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423553a8,
    48'h0000042355388,
    48'h000004235538c,
    48'h0000042355380,
    48'h0000042355384,
    48'h0000042355390,
    48'h0000042355378,
    48'h0000042355388,
    48'h0000042355388,
    48'h0000042355390,
    48'h0000042355378,
    48'h0000042355388,
    48'h000004214c8a8,
    48'h00000423553ac,
    48'h00000423553ac,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h00000423553ac,
    48'h00000423553a8,
    48'h00000423553ac,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h000004235538c,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042355390,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042355380,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042355384,
    48'h00000401367d0,
    48'h000007b0345c8,
    48'h0000040136428,
    48'h000007b034a48,
    48'h000004013893c,
    48'h0000042355378,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h000004235537a,
    48'h000004235537c,
    48'h0000042355368,
    48'h0000042355368,
    48'h0000042355368,
    48'h0000042355368,
    48'h0000042355368,
    48'h000004235536c,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042355370,
    48'h0000042355360,
    48'h0000042355364,
    48'h0000042355368,
    48'h0000042355370,
    48'h0000042355360,
    48'h000004235536c,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h0000042355390,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355380,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042355380,
    48'h0000042355384,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042355380,
    48'h0000040138938,
    48'h0000042355382,
    48'h000007b034f58,
    48'h0000042355384,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042355378,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042355378,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042355378,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042355378,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000000df84e8,
    48'h0000042355378,
    48'h0000000df84e9,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h000004235538c,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042355390,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042355380,
    48'h0000042355380,
    48'h0000042355384,
    48'h0000042355380,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000042355378,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000042355378,
    48'h000004235537a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042355390,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042355390,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034bac,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h00000423553a8,
    48'h0000042355388,
    48'h000004235538c,
    48'h0000042355380,
    48'h0000042355380,
    48'h0000042355380,
    48'h0000042355384,
    48'h0000042355382,
    48'h0000040001fac,
    48'h0000040023a68,
    48'h0000040023768,
    48'h000007b034e30,
    48'h0000040023760,
    48'h000007b034cc8,
    48'h00000423553b4,
    48'h0000042355398,
    48'h0000042355398,
    48'h000004213c310,
    48'h00000423553fc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af26c,
    48'h00000423553f0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423553f2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355400,
    48'h00000423553e0,
    48'h00000423553e4,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h000004235540c,
    48'h00000423b0422,
    48'h00000423b0428,
    48'h00000423553f0,
    48'h00000423553f0,
    48'h000004213c310,
    48'h000004235546c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af26c,
    48'h0000042355460,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355462,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355470,
    48'h0000042355450,
    48'h0000042355454,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235547c,
    48'h0000042355460,
    48'h0000042355460,
    48'h000004213c310,
    48'h00000423554e4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af26c,
    48'h00000423554d8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423554da,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423554e8,
    48'h00000423554c8,
    48'h00000423554cc,
    48'h0000042351df0,
    48'h00000423554c8,
    48'h00000423554c8,
    48'h00000423554d0,
    48'h00000423554b8,
    48'h00000423554c8,
    48'h000004214c8a8,
    48'h00000423554ec,
    48'h00000423554ec,
    48'h000007b03508c,
    48'h0000000dfcf58,
    48'h000007b035094,
    48'h0000000df7bf8,
    48'h000007b035094,
    48'h00000423554ec,
    48'h00000423554e8,
    48'h00000423554ec,
    48'h00000400025e4,
    48'h00000423554d0,
    48'h0000040139dd0,
    48'h00000423554bc,
    48'h0000040138938,
    48'h00000423554d0,
    48'h0000040139dd4,
    48'h00000423554c0,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df88e0,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9d80,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df88e4,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9d84,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df8444,
    48'h0000000df8445,
    48'h0000000df8446,
    48'h0000000df8447,
    48'h0000000df8448,
    48'h0000000df8449,
    48'h0000000df844a,
    48'h0000000df844b,
    48'h0000000df844c,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df8450,
    48'h0000000df8451,
    48'h0000000df8452,
    48'h0000000df8453,
    48'h0000000df8454,
    48'h0000000df8455,
    48'h0000000df8456,
    48'h0000000df8457,
    48'h0000000df8458,
    48'h0000040138938,
    48'h00000423554a8,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df8444,
    48'h0000040138938,
    48'h0000040139dd0,
    48'h00000423554aa,
    48'h00000423554ac,
    48'h0000042355498,
    48'h0000042355498,
    48'h0000042355498,
    48'h0000042355498,
    48'h0000042355498,
    48'h000004235549c,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423554a0,
    48'h0000042355490,
    48'h0000042355494,
    48'h0000042355498,
    48'h00000423554a0,
    48'h0000042355490,
    48'h000004235549c,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd0,
    48'h00000423554bc,
    48'h0000040138938,
    48'h000007b035050,
    48'h000004013893c,
    48'h00000423554b0,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df8450,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423554a8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df8444,
    48'h0000000df8444,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h00000423554a8,
    48'h0000000df8445,
    48'h00000423554a8,
    48'h0000000df8446,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h0000000df8447,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h00000423554a8,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423554b0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8450,
    48'h0000000df8450,
    48'h000007b0350bc,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h0000000df8451,
    48'h000007b034f5c,
    48'h0000040139a98,
    48'h000007b034f5c,
    48'h00000423554b0,
    48'h0000000df8452,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423554b0,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423554a8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df8448,
    48'h0000000df8448,
    48'h000007b0350bc,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h0000000df8449,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h00000423554a8,
    48'h0000000df844a,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423554b0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8453,
    48'h0000000df8453,
    48'h00000423554b0,
    48'h00000423554b4,
    48'h0000000df8454,
    48'h00000423554b0,
    48'h0000000df8455,
    48'h000007b034f5c,
    48'h0000040139a98,
    48'h000007b034f5c,
    48'h00000423554b0,
    48'h0000000df8456,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423554b0,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423554a8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df844b,
    48'h0000000df844b,
    48'h00000423554a8,
    48'h000007b034f40,
    48'h00000423554ac,
    48'h0000042355498,
    48'h0000000df844c,
    48'h000007b034f28,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h000007b0350a4,
    48'h00000423554a8,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423554b0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8457,
    48'h0000000df8457,
    48'h00000423554b0,
    48'h0000000df8458,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h000007b0350a4,
    48'h00000423554b0,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b034fd4,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423554bc,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423554c0,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000004013893c,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h000004013893c,
    48'h00000423554b4,
    48'h000007b034fa4,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h000007b034fa0,
    48'h000007b035018,
    48'h000007b035018,
    48'h0000040138938,
    48'h000007b035018,
    48'h000007b034fa0,
    48'h000007b035154,
    48'h000007b035018,
    48'h000007b035068,
    48'h000007b035150,
    48'h000007b035018,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb17b,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd0,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554aa,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423554bc,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423554bc,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fb8,
    48'h000007b035001,
    48'h000007b034fd4,
    48'h000007b034fec,
    48'h000007b035009,
    48'h000007b034fec,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb17c,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b4,
    48'h0000040136800,
    48'h0000040139540,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040139540,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c494,
    48'h000004214c69c,
    48'h0000040139544,
    48'h000004214c344,
    48'h000004013885c,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136514,
    48'h000004214c781,
    48'h000004214c599,
    48'h00000423554c0,
    48'h0000040136800,
    48'h0000040138f44,
    48'h00000423554c0,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h0000040022cc4,
    48'h0000040022de8,
    48'h0000040022ccc,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000004214c69c,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8018,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034bad,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000007b034ff4,
    48'h000004214c344,
    48'h000004013885c,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c344,
    48'h0000040139544,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h0000040021af0,
    48'h0000040021af8,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h0000040138eb0,
    48'h0000040138eb1,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h000007b034f4a,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h000007b034f48,
    48'h000007b034f4b,
    48'h000007b034f49,
    48'h000007b034f4b,
    48'h000007b034f49,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h0000040138eb1,
    48'h0000040138eb0,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c344,
    48'h000004214c69c,
    48'h000004214c494,
    48'h000004013885c,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c781,
    48'h000004013997c,
    48'h000004214c494,
    48'h00000423554b0,
    48'h0000040138f44,
    48'h00000423554b0,
    48'h000004214c494,
    48'h000004013997c,
    48'h000004214c69c,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c494,
    48'h0000040139544,
    48'h000007b035194,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554e0,
    48'h0000042355460,
    48'h0000042355460,
    48'h0000042355468,
    48'h00000423553f0,
    48'h00000423553f0,
    48'h000007b035154,
    48'h00000423553f4,
    48'h000004213a120,
    48'h0000042355400,
    48'h00000423553e0,
    48'h00000423553e8,
    48'h00000423553d0,
    48'h00000423554b0,
    48'h00000423553f8,
    48'h0000042355398,
    48'h0000042355398,
    48'h000007b035154,
    48'h000004235539c,
    48'h000004213a120,
    48'h00000423553a8,
    48'h0000042355388,
    48'h0000042355390,
    48'h0000042355378,
    48'h00000423554b0,
    48'h00000423553a0,
    48'h00000423550f8,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040139544,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040023890,
    48'h0000040023b38,
    48'h000007b034f11,
    48'h0000040139544,
    48'h0000040023b38,
    48'h0000040002490,
    48'h0000040023b38,
    48'h0000040001fac,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040001fac,
    48'h0000040023b38,
    48'h000007b034f11,
    48'h0000040023b38,
    48'h0000040023a5a,
    48'h00000400237b0,
    48'h0000040023898,
    48'h00000423b09e2,
    48'h000004013997c,
    48'h000007b034ff4,
    48'h000004013997c,
    48'h00000423b09e4,
    48'h00000401364c8,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c780,
    48'h0000040139978,
    48'h000004214c490,
    48'h00000423554a8,
    48'h0000040138f40,
    48'h00000423554a8,
    48'h000004214c490,
    48'h0000040139978,
    48'h000004214c698,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c490,
    48'h0000040139540,
    48'h000007b035194,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554ac,
    48'h00000423554a8,
    48'h0000042355498,
    48'h00000400015bc,
    48'h00000423554e0,
    48'h0000042355460,
    48'h0000042355460,
    48'h0000042355468,
    48'h00000423553f0,
    48'h00000423553f0,
    48'h000007b035154,
    48'h00000423553f4,
    48'h000004213a120,
    48'h0000042355400,
    48'h00000423553e0,
    48'h00000423553e4,
    48'h0000042351df0,
    48'h00000423553e8,
    48'h00000423553d0,
    48'h00000423553f8,
    48'h0000042355398,
    48'h0000042355398,
    48'h000007b035154,
    48'h000004235539c,
    48'h000004213a120,
    48'h00000423553a8,
    48'h0000042355388,
    48'h000004235538c,
    48'h0000042355380,
    48'h0000042355390,
    48'h00000423554a8,
    48'h0000042355378,
    48'h00000423554aa,
    48'h000004235537a,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h00000423554ac,
    48'h000004235537c,
    48'h0000042355498,
    48'h0000042355368,
    48'h000004235549a,
    48'h000004235536a,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h00000423554a0,
    48'h0000042355370,
    48'h0000042355490,
    48'h0000042355360,
    48'h0000042355494,
    48'h0000042355364,
    48'h0000042355390,
    48'h0000042355378,
    48'h00000423553a0,
    48'h00000423550f8,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff4,
    48'h000004013997c,
    48'h000004214c69c,
    48'h000004214c494,
    48'h00000423554b0,
    48'h0000040138f44,
    48'h00000423554b0,
    48'h00000400237b0,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000007b034fb8,
    48'h0000040139978,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h000004214c494,
    48'h000007b034fb9,
    48'h000004013997c,
    48'h00000423554b2,
    48'h000004214c344,
    48'h000004214c781,
    48'h00000423554b0,
    48'h00000423b09e2,
    48'h00000423554b0,
    48'h00000423554b2,
    48'h00000423554b0,
    48'h00000400015a4,
    48'h00000423554b0,
    48'h00000423b09e2,
    48'h000004213a240,
    48'h000004235914c,
    48'h0000000df7828,
    48'h000007b035258,
    48'h000007b03525c,
    48'h000007b035260,
    48'h000007b035264,
    48'h000007b035264,
    48'h000007b035260,
    48'h000004214c93c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b0a18,
    48'h00000423b0a18,
    48'h00000423b0a1a,
    48'h00000400020e0,
    48'h000004214c93c,
    48'h00000003840fc,
    48'h000007b03525c,
    48'h00000423b0a1c,
    48'h000004214c93c,
    48'h00000003840fd,
    48'h000007b035258,
    48'h00000423b0a20,
    48'h000004214c93c,
    48'h00000423b0a18,
    48'h000004214c90c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b0a28,
    48'h00000423b0a28,
    48'h00000423b0a3c,
    48'h00000423b0a40,
    48'h00000423b0a38,
    48'h00000423b0a44,
    48'h0000040002394,
    48'h0000040002394,
    48'h00000423b0a2c,
    48'h00000423554e0,
    48'h00000423b0a34,
    48'h00000423b0a30,
    48'h00000423b0a30,
    48'h000004235546c,
    48'h00000423554e0,
    48'h00000400015a4,
    48'h000007b034fb9,
    48'h000004214c69c,
    48'h000007b034ff4,
    48'h0000040023978,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h000004013997c,
    48'h00000423b09e2,
    48'h0000040022ccc,
    48'h0000040022cc4,
    48'h00000423554c0,
    48'h0000040022de8,
    48'h00000423554e8,
    48'h00000423554c8,
    48'h00000423554cc,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h00000423554f4,
    48'h00000423554d8,
    48'h00000423554d8,
    48'h000004213c310,
    48'h0000042355554,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af270,
    48'h0000042355548,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235554a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355558,
    48'h0000042355538,
    48'h000004235553c,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042355564,
    48'h0000042355548,
    48'h0000042355548,
    48'h000004213c310,
    48'h000004235534c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af270,
    48'h0000042355340,
    48'h0000042355340,
    48'h0000042355340,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042355340,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423555e4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h00000423555d8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423555da,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423555e8,
    48'h00000423555c8,
    48'h00000423555cc,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h0000042354c72,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h0000040023760,
    48'h000007b034ca8,
    48'h00000423555f4,
    48'h00000423555d8,
    48'h00000423555d8,
    48'h000004213c310,
    48'h000004235560c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042355600,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355602,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355610,
    48'h00000423555f8,
    48'h00000423555f8,
    48'h000004235561c,
    48'h00000423b0442,
    48'h00000423b0448,
    48'h0000042355600,
    48'h0000042355600,
    48'h000004213c310,
    48'h000004235564c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042355640,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355642,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355650,
    48'h0000042355630,
    48'h0000042355634,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235565c,
    48'h0000042355640,
    48'h0000042355640,
    48'h000004213c310,
    48'h0000042355674,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042355668,
    48'h0000042355668,
    48'h0000042355668,
    48'h0000042355668,
    48'h000004213c310,
    48'h0000042355684,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042355678,
    48'h0000042355678,
    48'h0000042355678,
    48'h0000042355678,
    48'h000004213c310,
    48'h0000042354f84,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042354f78,
    48'h0000042354f78,
    48'h0000042354f78,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042354f78,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423556d4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h00000423556c8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423556ca,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423556d8,
    48'h00000423556b8,
    48'h00000423556bc,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000423556c0,
    48'h00000423556b0,
    48'h00000423556b8,
    48'h00000423556b8,
    48'h00000423556c0,
    48'h00000423556b0,
    48'h00000423556b8,
    48'h000004214c8a8,
    48'h00000423556dc,
    48'h00000423556dc,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h00000423556dc,
    48'h00000423556d8,
    48'h00000423556dc,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423556bc,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423556c0,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354d00,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040136428,
    48'h000007b034a54,
    48'h000004013893c,
    48'h00000423556b0,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423556b2,
    48'h00000423556b4,
    48'h00000423556a0,
    48'h00000423556a0,
    48'h00000423556a0,
    48'h00000423556a0,
    48'h00000423556a0,
    48'h00000423556a4,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000423556a8,
    48'h0000042355698,
    48'h000004235569c,
    48'h00000423556a0,
    48'h00000423556a8,
    48'h0000042355698,
    48'h00000423556a4,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040139dd4,
    48'h00000423556c0,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042354d00,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042354d00,
    48'h0000040138938,
    48'h0000042354d02,
    48'h000007b034f58,
    48'h0000042354d04,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423556b0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h00000423556b0,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h00000423556b0,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h00000423556b0,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h0000000df84e8,
    48'h00000423556b0,
    48'h0000000df84e9,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423556bc,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423556c0,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042354d00,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423556c0,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423556c0,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034baf,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h00000423556d8,
    48'h00000423556b8,
    48'h00000423556bc,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042354d02,
    48'h0000040001fac,
    48'h0000040023a6e,
    48'h0000040023768,
    48'h000007b034e33,
    48'h0000040023760,
    48'h000007b034cd4,
    48'h00000423556e4,
    48'h00000423556c8,
    48'h00000423556c8,
    48'h000004213c310,
    48'h000004235572c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042355720,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355722,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h0000042355730,
    48'h0000042355710,
    48'h0000042355714,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042355718,
    48'h0000042355708,
    48'h0000042355710,
    48'h0000042355710,
    48'h0000042355718,
    48'h0000042355708,
    48'h0000042355710,
    48'h000004214c8a8,
    48'h0000042355734,
    48'h0000042355734,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h0000042355734,
    48'h0000042355730,
    48'h0000042355734,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h0000042355714,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042355718,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040136428,
    48'h000007b034a50,
    48'h000004013893c,
    48'h0000042355708,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h000004235570a,
    48'h000004235570c,
    48'h00000423556f8,
    48'h00000423556f8,
    48'h00000423556f8,
    48'h00000423556f8,
    48'h00000423556f8,
    48'h00000423556fc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042355700,
    48'h00000423556f0,
    48'h00000423556f4,
    48'h00000423556f8,
    48'h0000042355700,
    48'h00000423556f0,
    48'h00000423556fc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h0000042355718,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042354d90,
    48'h0000040138938,
    48'h0000042354d92,
    48'h000007b034f58,
    48'h0000042354d94,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042355708,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042355708,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042355708,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042355708,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000000df84e8,
    48'h0000042355708,
    48'h0000000df84e9,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h0000042355714,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042355718,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d90,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000042355708,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000042355708,
    48'h000004235570a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042355718,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042355718,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034baf,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000042355730,
    48'h0000042355710,
    48'h0000042355714,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d92,
    48'h0000040001fac,
    48'h0000040023a6c,
    48'h0000040023768,
    48'h000007b034e32,
    48'h0000040023760,
    48'h000007b034cd0,
    48'h000004235573c,
    48'h0000042355720,
    48'h0000042355720,
    48'h000004213c310,
    48'h0000042355784,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042355778,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235577a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355788,
    48'h0000042355750,
    48'h0000042355754,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h0000040023a5e,
    48'h0000040023768,
    48'h000007b034e2b,
    48'h0000040023760,
    48'h000007b034cb4,
    48'h0000042355794,
    48'h0000042355778,
    48'h0000042355778,
    48'h000004213c310,
    48'h0000042354fac,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042354fa0,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354fa2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042354fb0,
    48'h0000042354f90,
    48'h0000042354f94,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042354fbc,
    48'h0000042354fa0,
    48'h0000042354fa0,
    48'h000004213c310,
    48'h000004235501c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042355010,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355012,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355020,
    48'h0000042355000,
    48'h0000042355004,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235502c,
    48'h0000042355010,
    48'h0000042355010,
    48'h000004213c310,
    48'h000004235586c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042355860,
    48'h0000042355860,
    48'h0000042355860,
    48'h0000042355860,
    48'h000004213c310,
    48'h00000423b034c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h00000423b0340,
    48'h00000423b0340,
    48'h00000423b0340,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h00000423b0340,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h0000042354f54,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af27c,
    48'h0000042354f48,
    48'h0000042354f48,
    48'h0000042354f48,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042354f48,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423558c4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af280,
    48'h00000423558b8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423558ba,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423558c8,
    48'h00000423558a8,
    48'h00000423558ac,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h00000423558d4,
    48'h00000423b0462,
    48'h00000423b0468,
    48'h00000423558b8,
    48'h00000423558b8,
    48'h000004213c310,
    48'h0000042355934,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af280,
    48'h0000042355928,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235592a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355938,
    48'h0000042355918,
    48'h000004235591c,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042355944,
    48'h0000042355928,
    48'h0000042355928,
    48'h000004213c310,
    48'h000004235596c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af280,
    48'h0000042355960,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355962,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355970,
    48'h0000042355950,
    48'h0000042355954,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h000004235597c,
    48'h00000423b0472,
    48'h00000423b0478,
    48'h0000042355960,
    48'h0000042355960,
    48'h000004213c310,
    48'h00000423559dc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af284,
    48'h00000423559d0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423559d2,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423559e0,
    48'h00000423559c0,
    48'h00000423559c4,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h00000423559ec,
    48'h00000423559d0,
    48'h00000423559d0,
    48'h000004213c310,
    48'h000004235589c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af284,
    48'h0000042355890,
    48'h0000042355890,
    48'h0000042355890,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042355890,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423acd0c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h00000423acd00,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acd02,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423acd10,
    48'h00000423accf0,
    48'h00000423accf4,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h0000042354c72,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h0000040023760,
    48'h000007b034ca8,
    48'h00000423acd1c,
    48'h00000423acd00,
    48'h00000423acd00,
    48'h000004213c310,
    48'h00000423acd34,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h00000423acd28,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acd2a,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423acd38,
    48'h00000423acd20,
    48'h00000423acd20,
    48'h00000423acd44,
    48'h00000423b0482,
    48'h00000423b0488,
    48'h00000423acd28,
    48'h00000423acd28,
    48'h000004213c310,
    48'h00000423acd74,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h00000423acd68,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acd6a,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423acd78,
    48'h00000423acd58,
    48'h00000423acd5c,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h00000423acd84,
    48'h00000423acd68,
    48'h00000423acd68,
    48'h000004213c310,
    48'h00000423acd9c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h00000423acd90,
    48'h00000423acd90,
    48'h00000423acd90,
    48'h00000423acd90,
    48'h000004213c310,
    48'h0000042355884,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h0000042355878,
    48'h0000042355878,
    48'h0000042355878,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042355878,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423acde4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423acdd8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acdda,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423acde8,
    48'h00000423acdc8,
    48'h00000423acdcc,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h00000423acdd0,
    48'h00000423acdb8,
    48'h00000423acdc8,
    48'h00000423acdc8,
    48'h00000423acdd0,
    48'h00000423acdb8,
    48'h00000423acdc8,
    48'h000004214c8a8,
    48'h00000423acdec,
    48'h00000423acdec,
    48'h000007b03508c,
    48'h0000000dfd1c8,
    48'h000007b035094,
    48'h0000000df7e68,
    48'h000007b035094,
    48'h00000423acdec,
    48'h00000423acde8,
    48'h00000423acdec,
    48'h0000040002854,
    48'h0000040139dd0,
    48'h00000423acdcc,
    48'h0000040138938,
    48'h00000423acdd0,
    48'h0000040139dd4,
    48'h00000423acdbc,
    48'h000004013893c,
    48'h00000423acdd0,
    48'h0000040139dd8,
    48'h00000423acdc0,
    48'h0000040138940,
    48'h000007b03508c,
    48'h0000000df9510,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000dfa9b0,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df9514,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000dfa9b4,
    48'h000007b03506c,
    48'h000007b03508c,
    48'h0000000df9518,
    48'h000007b034f18,
    48'h000007b034f30,
    48'h0000000dfa9b8,
    48'h000007b035070,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df85f0,
    48'h0000000df85f1,
    48'h0000000df85f2,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df85f4,
    48'h0000040138938,
    48'h000004013893c,
    48'h00000423acdb0,
    48'h0000042354e20,
    48'h00000423acdb4,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h000007b035031,
    48'h0000000df85f5,
    48'h0000040138940,
    48'h000007b035058,
    48'h000007b034f30,
    48'h0000000df8750,
    48'h0000000df8751,
    48'h0000000df8752,
    48'h0000040138938,
    48'h00000423acdb0,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df85f0,
    48'h0000040138938,
    48'h00000423acdb4,
    48'h00000401367d0,
    48'h000007b0345a8,
    48'h0000040136428,
    48'h000007b034a28,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df85f4,
    48'h000004013893c,
    48'h0000042354e24,
    48'h00000401367d0,
    48'h000007b0345b4,
    48'h0000040136428,
    48'h000007b034a34,
    48'h0000040138940,
    48'h00000423acda8,
    48'h000007b035020,
    48'h000007b034f48,
    48'h000007b034f30,
    48'h0000000df8750,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acdb0,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df85f0,
    48'h0000000df85f0,
    48'h000007b035018,
    48'h0000000df85f1,
    48'h000007b034f58,
    48'h0000040139a84,
    48'h000007b034f58,
    48'h00000423acdb0,
    48'h0000040138938,
    48'h00000423acdb2,
    48'h000007b034f58,
    48'h00000423acdb4,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df85f2,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df85f4,
    48'h0000000df85f4,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035031,
    48'h000007b034f70,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b034f58,
    48'h000007b035150,
    48'h000007b035154,
    48'h000004013893c,
    48'h0000040138938,
    48'h0000040139dd4,
    48'h0000040139dd0,
    48'h000007b035154,
    48'h000007b035150,
    48'h00000423acdb0,
    48'h0000042354e20,
    48'h00000423acdb2,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h0000040001fac,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h0000040139db0,
    48'h00000423acdbc,
    48'h0000040138950,
    48'h00000423afb50,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h0000040022e60,
    48'h00000423acde8,
    48'h00000423acdc8,
    48'h00000423acdcc,
    48'h00000423acdb0,
    48'h00000423acdd0,
    48'h00000423acdb8,
    48'h000004214c9c0,
    48'h0000040002164,
    48'h00000003840fd,
    48'h00000423acdc0,
    48'h00000423acda8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h00000003840fc,
    48'h00000423acdbc,
    48'h0000042351df8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h0000040002490,
    48'h00000423acdbc,
    48'h0000040022e70,
    48'h0000042354e20,
    48'h0000040022e60,
    48'h00000423acdb4,
    48'h00000423acdf4,
    48'h00000423b0522,
    48'h00000423b0524,
    48'h0000042354e24,
    48'h00000423b0528,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df85f5,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h0000042354e20,
    48'h000007b034f5c,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423acda8,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df8750,
    48'h0000000df8750,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423acda8,
    48'h0000000df8751,
    48'h00000423acda8,
    48'h00000423acdac,
    48'h0000000df8752,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b0350bc,
    48'h000007b034f72,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b034f60,
    48'h000007b034fa8,
    48'h000007b034f72,
    48'h000007b035002,
    48'h000007b034f7a,
    48'h000007b03500a,
    48'h000007b034f90,
    48'h000007b034fd8,
    48'h000007b034f82,
    48'h000007b035012,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b034ff0,
    48'h000007b035000,
    48'h000007b034fd0,
    48'h000007b035001,
    48'h000007b034fd4,
    48'h000007b034fe8,
    48'h000007b035002,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423acdcc,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423acdbc,
    48'h000007b034fbc,
    48'h0000040139dd8,
    48'h000007b035058,
    48'h00000423acdc0,
    48'h000007b034fc0,
    48'h000007b035000,
    48'h0000040138938,
    48'h00000423acdb0,
    48'h00000423acdb0,
    48'h000007b035001,
    48'h000004013893c,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h000007b035002,
    48'h000007b035000,
    48'h000007b034fd0,
    48'h000007b034fe8,
    48'h000007b035018,
    48'h000007b035018,
    48'h000007b034fe8,
    48'h000007b03501c,
    48'h000007b034fa0,
    48'h000007b035154,
    48'h000007b034fe8,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b035068,
    48'h000007b035148,
    48'h000007b035144,
    48'h000007b03514c,
    48'h000004013893c,
    48'h0000040138938,
    48'h0000040139dd4,
    48'h0000040139dd0,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h0000042354e20,
    48'h0000042354e22,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423acdbc,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423acdbc,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h0000040022cc4,
    48'h0000040022de8,
    48'h0000040022ccc,
    48'h0000040139978,
    48'h0000040139540,
    48'h000007b035210,
    48'h000007b035214,
    48'h000007b035214,
    48'h000007b035210,
    48'h00000423acdb0,
    48'h0000042354e20,
    48'h00000423acdb2,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h0000040001fac,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h0000040139db0,
    48'h00000423acdbc,
    48'h0000040138950,
    48'h00000423afb50,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h0000040022e60,
    48'h00000423acde8,
    48'h00000423acdc8,
    48'h00000423acdcc,
    48'h00000423acdb0,
    48'h00000423acdd0,
    48'h00000423acdb8,
    48'h000004214c9c0,
    48'h0000040002164,
    48'h00000003840fd,
    48'h00000423acdc0,
    48'h00000423acda8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h00000003840fc,
    48'h00000423acdbc,
    48'h0000042351df8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h0000040002490,
    48'h00000423acdbc,
    48'h0000040022e70,
    48'h0000042354e20,
    48'h0000040022e60,
    48'h00000423acdb4,
    48'h00000423acdf4,
    48'h00000423b0522,
    48'h00000423b0524,
    48'h0000042354e24,
    48'h00000423b0528,
    48'h0000040139978,
    48'h0000042354e20,
    48'h000007b03520c,
    48'h000007b035210,
    48'h0000040022e78,
    48'h000007b035214,
    48'h0000040022e60,
    48'h00000423acdb4,
    48'h000007b035254,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423acde0,
    48'h0000042355878,
    48'h0000040022e88,
    48'h000007b034fe8,
    48'h000007b034fbc,
    48'h0000040022e88,
    48'h000007b034fb8,
    48'h000007b035001,
    48'h000007b034fd4,
    48'h000007b035002,
    48'h000007b034ff0,
    48'h000007b034fd8,
    48'h00000400015a4,
    48'h0000040138940,
    48'h00000423acda8,
    48'h00000423acda8,
    48'h00000423acda8,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040138eb0,
    48'h000004214c490,
    48'h000007b03508c,
    48'h0000000df8288,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034bb4,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001fac,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h0000040138858,
    48'h0000040001fac,
    48'h0000040001fac,
    48'h000004214c780,
    48'h0000040139978,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h0000040023760,
    48'h0000040023768,
    48'h000007b034ca8,
    48'h000007b034e28,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000007b034fb8,
    48'h0000040139978,
    48'h0000042354e22,
    48'h000004214c780,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423acdb2,
    48'h0000042354e20,
    48'h0000042354e22,
    48'h0000042354e20,
    48'h00000400015a4,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423acdb2,
    48'h000004213a240,
    48'h000004235914c,
    48'h0000000df7828,
    48'h000007b035258,
    48'h000007b03525c,
    48'h000007b035260,
    48'h000007b035264,
    48'h000007b035264,
    48'h000007b035260,
    48'h000004214c93c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b0a48,
    48'h00000423b0a48,
    48'h00000423b0a4a,
    48'h00000400020e0,
    48'h000004214c93c,
    48'h00000003840fc,
    48'h000007b03525c,
    48'h00000423b0a4c,
    48'h000004214c93c,
    48'h00000003840fd,
    48'h000007b035258,
    48'h00000423b0a50,
    48'h000004214c93c,
    48'h00000423b0a48,
    48'h000004214c90c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b0a58,
    48'h00000423b0a58,
    48'h00000423b0a6c,
    48'h00000423b0a70,
    48'h00000423b0a68,
    48'h00000423b0a74,
    48'h0000040002394,
    48'h0000040002394,
    48'h00000423b0a5c,
    48'h00000423acde0,
    48'h00000423b0a64,
    48'h00000423b0a60,
    48'h00000423b0a60,
    48'h0000042355884,
    48'h00000423acde0,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h0000040139978,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h00000423acdb2,
    48'h0000040022cc0,
    48'h0000040022cb8,
    48'h00000423acdbc,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h0000040139978,
    48'h00000423acdb2,
    48'h0000040022ccc,
    48'h0000040022cc4,
    48'h00000423acdcc,
    48'h0000040022de8,
    48'h00000423acde8,
    48'h00000423acdc8,
    48'h00000423acdcc,
    48'h00000423acdb0,
    48'h00000423acdb0,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h00000423acdf4,
    48'h00000423b0522,
    48'h00000423b0528,
    48'h00000423acdd8,
    48'h00000423acdd8,
    48'h000004213c310,
    48'h00000423ace24,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423ace18,
    48'h00000423ace18,
    48'h00000423ace18,
    48'h00000423ace18,
    48'h000004213c310,
    48'h00000423ace6c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423ace60,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423ace62,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423ace70,
    48'h00000423ace50,
    48'h00000423ace54,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h00000423ace3c,
    48'h00000423ace3a,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h0000040023760,
    48'h000007b034ca8,
    48'h00000423ace7c,
    48'h00000423b0502,
    48'h00000423b0508,
    48'h00000423ace60,
    48'h00000423ace60,
    48'h000004213c310,
    48'h00000423aceac,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423acea0,
    48'h00000423acea0,
    48'h00000423acea0,
    48'h00000423acea0,
    48'h000004213c310,
    48'h00000423acefc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423acef0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acef2,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423acf00,
    48'h00000423acee0,
    48'h00000423acee4,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h00000423acee8,
    48'h00000423b0860,
    48'h00000423acee0,
    48'h00000423acee0,
    48'h00000423acee8,
    48'h00000423b0860,
    48'h00000423acee0,
    48'h000004214c8a8,
    48'h00000423acf04,
    48'h00000423acf04,
    48'h000007b03508c,
    48'h0000000dfd13c,
    48'h000007b035094,
    48'h0000000df7ddc,
    48'h000007b035094,
    48'h00000423acf04,
    48'h00000423acf00,
    48'h00000423acf04,
    48'h00000400027c8,
    48'h0000040139dd0,
    48'h00000423acee4,
    48'h0000040138938,
    48'h00000423acee8,
    48'h0000040139dd4,
    48'h00000423b0864,
    48'h000004013893c,
    48'h00000423acee8,
    48'h0000040139dd8,
    48'h00000423b0868,
    48'h0000040138940,
    48'h000007b03508c,
    48'h0000000df9254,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000dfa6f4,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df9258,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000dfa6f8,
    48'h000007b03506c,
    48'h000007b03508c,
    48'h0000000df925c,
    48'h000007b034f18,
    48'h000007b034f30,
    48'h0000000dfa6fc,
    48'h000007b035070,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df868c,
    48'h0000000df868d,
    48'h0000000df868e,
    48'h0000000df868f,
    48'h0000000df8690,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df8674,
    48'h0000000df8675,
    48'h0000040138938,
    48'h000004013893c,
    48'h00000423acec8,
    48'h00000423ace38,
    48'h00000423acecc,
    48'h00000423ace38,
    48'h00000423ace3c,
    48'h000007b035031,
    48'h0000040138938,
    48'h0000040138940,
    48'h00000423acec8,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h000007b035032,
    48'h0000000df8676,
    48'h0000000df8677,
    48'h0000040138938,
    48'h000004013893c,
    48'h00000423acec8,
    48'h00000423ace38,
    48'h00000423acecc,
    48'h00000423ace38,
    48'h00000423ace3c,
    48'h000007b035031,
    48'h0000040138938,
    48'h0000040138940,
    48'h00000423acec8,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h000007b035032,
    48'h0000000df8678,
    48'h0000040138940,
    48'h000007b035058,
    48'h000007b034f30,
    48'h0000000df8728,
    48'h0000000df8729,
    48'h0000000df872a,
    48'h0000000df872b,
    48'h0000000df872c,
    48'h0000000df872d,
    48'h0000000df872e,
    48'h0000000df872f,
    48'h0000000df8730,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df868c,
    48'h0000040138938,
    48'h00000423acecc,
    48'h00000401367d0,
    48'h000007b0345a8,
    48'h0000040136428,
    48'h000007b034a28,
    48'h000004013893c,
    48'h00000423ace38,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df8674,
    48'h000004013893c,
    48'h00000423ace3c,
    48'h00000401367d0,
    48'h000007b0345a8,
    48'h0000040136428,
    48'h000007b034a28,
    48'h0000040138940,
    48'h00000423b0848,
    48'h000007b035020,
    48'h000007b034f48,
    48'h000007b034f30,
    48'h0000000df8728,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df868c,
    48'h0000000df868c,
    48'h000007b035018,
    48'h0000000df868d,
    48'h000007b0350bc,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h00000423acec8,
    48'h00000423acec8,
    48'h0000000df868e,
    48'h000007b034f28,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h000007b0350a4,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f88,
    48'h000007b0350a4,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423ace38,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8674,
    48'h0000000df8674,
    48'h0000000df8675,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035031,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df8676,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423ace38,
    48'h000007b034f5c,
    48'h000007b034f8c,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423b0848,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df8728,
    48'h0000000df8728,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423b0848,
    48'h0000000df8729,
    48'h00000423b0848,
    48'h00000423b084c,
    48'h0000000df872a,
    48'h00000423b0848,
    48'h0000000df872b,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b034f7a,
    48'h00000423b0848,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df868f,
    48'h0000000df868f,
    48'h000007b034f58,
    48'h0000040139a84,
    48'h000007b034f58,
    48'h00000423acec8,
    48'h0000040138938,
    48'h00000423aceca,
    48'h000007b034f58,
    48'h00000423acecc,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df8690,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423ace38,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8677,
    48'h0000000df8677,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035031,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df8678,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423b0848,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df872c,
    48'h0000000df872c,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423b0848,
    48'h0000000df872d,
    48'h000007b0350bc,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h0000000df872e,
    48'h00000423b0848,
    48'h00000423b084c,
    48'h0000000df872f,
    48'h00000423b0848,
    48'h0000000df8730,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b034f7a,
    48'h00000423b0848,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b034f60,
    48'h000007b034fa8,
    48'h000007b034f72,
    48'h000007b035002,
    48'h000007b034f7a,
    48'h000007b03500a,
    48'h000007b034f90,
    48'h000007b034fd8,
    48'h000007b034f82,
    48'h000007b035012,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b03509c,
    48'h000007b03509c,
    48'h000007b035058,
    48'h000004013893c,
    48'h000007b035054,
    48'h0000040138940,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df868c,
    48'h0000000df868c,
    48'h000007b035018,
    48'h0000000df868d,
    48'h000007b0350bc,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h00000423acec8,
    48'h00000423acec8,
    48'h0000000df868e,
    48'h000007b034f28,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h000007b0350a4,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f88,
    48'h000007b0350a4,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423b0848,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8674,
    48'h0000000df8674,
    48'h0000000df8675,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035032,
    48'h000007b034f70,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b035150,
    48'h000007b035154,
    48'h000004013893c,
    48'h0000040138938,
    48'h0000040139dd4,
    48'h0000040139dd0,
    48'h000007b035154,
    48'h000007b035150,
    48'h00000423acec8,
    48'h00000423b0848,
    48'h00000423aceca,
    48'h00000423b084a,
    48'h0000040001fac,
    48'h0000040001f9c,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h0000040139db0,
    48'h00000423b0864,
    48'h0000040138950,
    48'h00000423afb50,
    48'h00000423aceca,
    48'h0000040001fac,
    48'h0000040022e60,
    48'h00000423acf00,
    48'h00000423acee0,
    48'h00000423acee4,
    48'h00000423acec8,
    48'h00000423acee8,
    48'h00000423b0860,
    48'h000004214c9ac,
    48'h0000040002150,
    48'h00000003840fd,
    48'h00000423b0868,
    48'h00000423b0848,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h00000003840fc,
    48'h00000423b0864,
    48'h0000042351df8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h0000040002468,
    48'h00000423b0864,
    48'h0000040022e70,
    48'h00000423b0848,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df8676,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423b0848,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423ace38,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df8728,
    48'h0000000df8728,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423ace38,
    48'h0000040138940,
    48'h00000423ace3a,
    48'h000007b034f60,
    48'h00000423ace3c,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df8729,
    48'h00000423ace38,
    48'h0000000df872a,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h0000000df872b,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b0350bc,
    48'h000007b034f72,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df868f,
    48'h0000000df868f,
    48'h000007b034f58,
    48'h0000040139a84,
    48'h000007b034f58,
    48'h00000423acec8,
    48'h0000040138938,
    48'h00000423aceca,
    48'h000007b034f58,
    48'h00000423acecc,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df8690,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423b0848,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8677,
    48'h0000000df8677,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035032,
    48'h000007b034f70,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b034f58,
    48'h000007b035150,
    48'h000007b035154,
    48'h000004013893c,
    48'h0000040138938,
    48'h0000040139dd4,
    48'h0000040139dd0,
    48'h000007b035154,
    48'h000007b035150,
    48'h00000423acec8,
    48'h00000423b0848,
    48'h00000423aceca,
    48'h00000423b084a,
    48'h0000040001fac,
    48'h0000040001f9c,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h0000040139db0,
    48'h00000423b0864,
    48'h0000040138950,
    48'h00000423afb50,
    48'h00000423aceca,
    48'h0000040001fac,
    48'h0000040022e60,
    48'h00000423acf00,
    48'h00000423acee0,
    48'h00000423acee4,
    48'h00000423acec8,
    48'h00000423acee8,
    48'h00000423b0860,
    48'h000004214c9ac,
    48'h0000040002150,
    48'h00000003840fd,
    48'h00000423b0868,
    48'h00000423b0848,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h00000003840fc,
    48'h00000423b0864,
    48'h0000042351df8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h0000040002490,
    48'h00000423b0864,
    48'h0000040022e70,
    48'h00000423b0848,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df8678,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423b0848,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423ace38,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df872c,
    48'h0000000df872c,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423ace38,
    48'h0000040138940,
    48'h00000423ace3a,
    48'h000007b034f60,
    48'h00000423ace3c,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df872d,
    48'h000007b0350bc,
    48'h00000423ace38,
    48'h00000423ace3c,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h0000000df872e,
    48'h00000423ace38,
    48'h0000000df872f,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h0000000df8730,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b0350bc,
    48'h000007b034f72,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b03509c,
    48'h000007b03509c,
    48'h000007b035054,
    48'h000004013893c,
    48'h000007b035058,
    48'h0000040138940,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b034ff0,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035002,
    48'h000007b034fd8,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423acee4,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423b0864,
    48'h000007b034fbc,
    48'h0000040139dd8,
    48'h000007b035058,
    48'h00000400341a0,
    48'h0000000dfcfa8,
    48'h000007b034dd4,
    48'h0000000df7c48,
    48'h000007b034dd4,
    48'h00000423aebbc,
    48'h00000423aebb8,
    48'h00000423aebbc,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423aeb9c,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423aeba0,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df8a70,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9f10,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8a74,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000df9f14,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h00000423aeb90,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000040139dd0,
    48'h00000423aeb92,
    48'h00000423aeb94,
    48'h00000423aeb88,
    48'h00000423aeb88,
    48'h00000423aeb88,
    48'h00000423aeb88,
    48'h00000423aeb8c,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h00000423aeb88,
    48'h0000040022e80,
    48'h00000423aeb88,
    48'h000004214c9d4,
    48'h0000040002178,
    48'h0000000384130,
    48'h00000423aeb8c,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h00000401367d0,
    48'h000007b0345e4,
    48'h00000423aeb8c,
    48'h00000423aeb94,
    48'h0000040022e80,
    48'h0000040139dd0,
    48'h00000423aeb9c,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000004013893c,
    48'h00000423aeb80,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423aeb82,
    48'h00000423aeb84,
    48'h00000423aeb70,
    48'h00000423aeb70,
    48'h00000423aeb70,
    48'h00000423aeb70,
    48'h00000423aeb70,
    48'h00000423aeb74,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423aeb78,
    48'h00000423aeb68,
    48'h00000423aeb6c,
    48'h00000423aeb70,
    48'h00000423aeb78,
    48'h00000423aeb68,
    48'h00000423aeb74,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h00000423aeba0,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h00000423aeb90,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b034d58,
    48'h0000000df84d5,
    48'h000007b034dfc,
    48'h00000423aeb90,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h00000423aeb90,
    48'h0000000df84d6,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h00000423aeb80,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034c9c,
    48'h0000040139a84,
    48'h000007b034c9c,
    48'h00000423aeb80,
    48'h0000000df84e5,
    48'h000007b034c9c,
    48'h0000040139bac,
    48'h000007b034c9c,
    48'h00000423aeb80,
    48'h0000000df84e6,
    48'h000007b034c9c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034c9c,
    48'h00000423aeb80,
    48'h0000000df84e7,
    48'h000007b034dfc,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h0000000df84e8,
    48'h00000423aeb80,
    48'h0000000df84e9,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h0000000df84ea,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423aeb9c,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423aeba0,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h00000423aeb90,
    48'h00000423aeb90,
    48'h00000423aeb90,
    48'h000007b034ce0,
    48'h000007b034d58,
    48'h00000423aeba8,
    48'h000007b034d58,
    48'h000007b034d58,
    48'h0000040138938,
    48'h000007b034ce0,
    48'h000007b034e94,
    48'h000007b034d58,
    48'h000007b034e90,
    48'h000007b034d58,
    48'h000007b034da8,
    48'h000007b034e8c,
    48'h000007b034dcc,
    48'h0000000dfb1df,
    48'h000007b034e88,
    48'h000007b034e84,
    48'h0000040139dd0,
    48'h000007b034e90,
    48'h000007b034e8c,
    48'h000007b034e88,
    48'h000007b034e94,
    48'h00000423aeb90,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423aeb9c,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000040022cb0,
    48'h0000040022e88,
    48'h000007b034cf8,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h000007b034ce4,
    48'h000007b034d5c,
    48'h000007b034d5c,
    48'h000004013893c,
    48'h000007b034d5c,
    48'h000007b034ce4,
    48'h000007b034e94,
    48'h000007b034d5c,
    48'h000007b034dac,
    48'h000007b034e90,
    48'h000007b034d5c,
    48'h000007b034e8c,
    48'h000007b034dcc,
    48'h0000000dfb1e0,
    48'h000007b034e88,
    48'h000007b034e84,
    48'h0000040139dd4,
    48'h000007b034e90,
    48'h000007b034e8c,
    48'h000007b034e88,
    48'h000007b034e94,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb80,
    48'h00000423aeb82,
    48'h0000040136800,
    48'h0000040139540,
    48'h000004214c780,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040139540,
    48'h000004214c780,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c494,
    48'h000004214c69c,
    48'h0000040139544,
    48'h000004214c344,
    48'h000004013885c,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136514,
    48'h000004214c781,
    48'h000004214c599,
    48'h00000423aeba0,
    48'h0000040136800,
    48'h0000040138f44,
    48'h00000423aeba0,
    48'h0000040022cb0,
    48'h000007b034cfc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000004214c69c,
    48'h0000040136800,
    48'h0000040138eb0,
    48'h000007b034dcc,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000007b03451c,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423aebaa,
    48'h000007b034390,
    48'h000007b0344a8,
    48'h000007b034400,
    48'h000007b0344e0,
    48'h000007b034394,
    48'h000007b0344ac,
    48'h000007b034404,
    48'h000007b0344e4,
    48'h000007b034398,
    48'h000007b0344b0,
    48'h000007b034408,
    48'h000007b0344e8,
    48'h000007b03439c,
    48'h000007b0344b4,
    48'h000007b03440c,
    48'h000007b0344ec,
    48'h000007b0343a0,
    48'h000007b0344b8,
    48'h000007b034410,
    48'h000007b0344f0,
    48'h000007b0343a4,
    48'h000007b0344bc,
    48'h000007b034414,
    48'h000007b0344f4,
    48'h000007b0343a8,
    48'h000007b0344c0,
    48'h000007b034418,
    48'h000007b0344f8,
    48'h000007b0343ac,
    48'h000007b0344c4,
    48'h000007b03441c,
    48'h000007b0344fc,
    48'h000007b0343b0,
    48'h000007b0344c8,
    48'h000007b034420,
    48'h000007b034500,
    48'h000007b0343b4,
    48'h000007b0344cc,
    48'h000007b034424,
    48'h000007b034504,
    48'h000007b0343b8,
    48'h000007b0344d0,
    48'h000007b034428,
    48'h000007b034508,
    48'h000007b0343bc,
    48'h000007b0344d4,
    48'h000007b03442c,
    48'h000007b03450c,
    48'h000007b0343c0,
    48'h000007b0344d8,
    48'h000007b034430,
    48'h000007b034510,
    48'h000007b0343c4,
    48'h000007b0344dc,
    48'h000007b034434,
    48'h000007b034514,
    48'h00000423aebb4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423aebe0,
    48'h00000423aebe0,
    48'h00000423aebec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423aec30,
    48'h00000423aec30,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423aec40,
    48'h00000423aec20,
    48'h000004214c8a8,
    48'h00000423aec44,
    48'h00000423aec44,
    48'h000007b034dcc,
    48'h0000000dfd2f8,
    48'h000007b034dd4,
    48'h0000000df7f98,
    48'h000007b034dd4,
    48'h00000423aec44,
    48'h00000423aec40,
    48'h00000423aec44,
    48'h0000040002984,
    48'h0000040139dd0,
    48'h00000423aec24,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423aec28,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df9b00,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000dfafa0,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df9b04,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000dfafa4,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df8778,
    48'h0000000df8779,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84f8,
    48'h0000000df84f9,
    48'h0000040138938,
    48'h00000423aec18,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df8778,
    48'h0000040138938,
    48'h0000040139dd0,
    48'h00000423aec1a,
    48'h00000423aec1c,
    48'h000004239fdc8,
    48'h000004239fdc8,
    48'h000004239fdc8,
    48'h0000040022e80,
    48'h000004239fdc8,
    48'h00000423aec1c,
    48'h0000040022e80,
    48'h0000040139dd0,
    48'h00000423aec24,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000004013893c,
    48'h00000423aec10,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84f8,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h00000423aec18,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df8778,
    48'h0000000df8778,
    48'h000007b034dfc,
    48'h00000423aec18,
    48'h00000423aec18,
    48'h00000423aec1a,
    48'h00000423aec1c,
    48'h000007b034f50,
    48'h000004239fdc8,
    48'h000004239fdc8,
    48'h00000423aec18,
    48'h00000423aec18,
    48'h000007b034df4,
    48'h0000000df8779,
    48'h000007b034c68,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h00000423aec10,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84f8,
    48'h0000000df84f8,
    48'h000007b034dfc,
    48'h00000423aec10,
    48'h000007b034c9c,
    48'h0000040139a98,
    48'h000007b034c9c,
    48'h00000423aec10,
    48'h0000000df84f9,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423aec24,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423aec28,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h00000423aec18,
    48'h00000423aec18,
    48'h00000423aec18,
    48'h000007b034ce0,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423aec10,
    48'h00000423aec10,
    48'h00000423aec10,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df83b8,
    48'h0000040136800,
    48'h00000423aec3c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423aec78,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423aec88,
    48'h00000423aec68,
    48'h00000423aec6c,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h00000423aec70,
    48'h00000423aec58,
    48'h00000423aec68,
    48'h00000423aec68,
    48'h00000423aec70,
    48'h00000423aec58,
    48'h00000423aec68,
    48'h000004214c8a8,
    48'h00000423aec8c,
    48'h00000423aec8c,
    48'h000007b034dcc,
    48'h0000000dfd064,
    48'h000007b034dd4,
    48'h0000000df7d04,
    48'h000007b034dd4,
    48'h00000423aec8c,
    48'h00000423aec88,
    48'h00000423aec8c,
    48'h00000400026f0,
    48'h0000040139dd0,
    48'h00000423aec6c,
    48'h0000040138938,
    48'h00000423aec70,
    48'h0000040139dd4,
    48'h00000423aec5c,
    48'h000004013893c,
    48'h00000423aec70,
    48'h0000040139dd8,
    48'h00000423aec60,
    48'h0000040138940,
    48'h000007b034dcc,
    48'h0000000df8e1c,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000dfa2bc,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8e20,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000dfa2c0,
    48'h000007b034dac,
    48'h000007b034dcc,
    48'h0000000df8e24,
    48'h000007b034c58,
    48'h000007b034c70,
    48'h0000000dfa2c4,
    48'h000007b034db0,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df863c,
    48'h0000000df863d,
    48'h0000000df863e,
    48'h0000000df863f,
    48'h0000000df8640,
    48'h0000000df8641,
    48'h0000000df8642,
    48'h0000000df8643,
    48'h0000000df8644,
    48'h0000000df8645,
    48'h0000000df8646,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df8648,
    48'h0000000df8649,
    48'h0000040138938,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034d71,
    48'h0000040138938,
    48'h0000040138940,
    48'h0000042351e38,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h000007b034d72,
    48'h0000000df864a,
    48'h0000000df864b,
    48'h0000040138938,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034d71,
    48'h0000040138938,
    48'h0000040138940,
    48'h0000042351e38,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h000007b034d72,
    48'h0000000df864c,
    48'h0000000df864d,
    48'h0000000df864e,
    48'h0000000df864f,
    48'h0000000df8650,
    48'h0000000df8651,
    48'h0000000df8652,
    48'h0000040138940,
    48'h000007b034d98,
    48'h000007b034c70,
    48'h0000000df8654,
    48'h0000000df8655,
    48'h0000000df8656,
    48'h0000000df8657,
    48'h0000000df8658,
    48'h0000000df8659,
    48'h0000000df865a,
    48'h0000000df865b,
    48'h0000000df865c,
    48'h0000000df865d,
    48'h0000000df865e,
    48'h0000000df865f,
    48'h0000000df8660,
    48'h0000000df8661,
    48'h0000000df8662,
    48'h0000000df8663,
    48'h0000000df8664,
    48'h0000000df8665,
    48'h0000000df8666,
    48'h0000040138938,
    48'h0000042351e38,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df863c,
    48'h0000040138938,
    48'h0000042351e3c,
    48'h00000401367d0,
    48'h000007b0345e4,
    48'h0000040136428,
    48'h000007b034a64,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df8648,
    48'h000004013893c,
    48'h0000042351e3c,
    48'h00000401367d0,
    48'h000007b0345e4,
    48'h0000040136428,
    48'h000007b034a64,
    48'h0000040138940,
    48'h00000423aec50,
    48'h000007b034d60,
    48'h000007b034c88,
    48'h000007b034c70,
    48'h0000000df8654,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042351e38,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df863c,
    48'h0000000df863c,
    48'h000007b034d58,
    48'h0000000df863d,
    48'h000007b034dfc,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h0000042351e38,
    48'h0000042351e38,
    48'h0000000df863e,
    48'h000007b034c68,
    48'h000007b034cc0,
    48'h000007b034cb8,
    48'h000007b034de4,
    48'h0000042351e38,
    48'h000007b034c98,
    48'h000007b034cc8,
    48'h000007b034de4,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df8648,
    48'h0000000df8648,
    48'h0000000df8649,
    48'h000007b034ccc,
    48'h000007b034ddc,
    48'h000007b034d71,
    48'h000007b034cb0,
    48'h000007b034c98,
    48'h000007b034c9c,
    48'h0000000df864a,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034cb9,
    48'h0000042351e38,
    48'h000007b034c9c,
    48'h000007b034ccc,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h00000423aec50,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df8654,
    48'h0000000df8654,
    48'h000007b034ca0,
    48'h0000040139a84,
    48'h000007b034ca0,
    48'h00000423aec50,
    48'h0000000df8655,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8656,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8657,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8658,
    48'h00000423aec50,
    48'h0000000df8659,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034cba,
    48'h00000423aec50,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034dec,
    48'h000007b034de4,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042351e38,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df863f,
    48'h0000000df863f,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042351e38,
    48'h0000040138938,
    48'h0000042351e3a,
    48'h000007b034c98,
    48'h0000042351e3c,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df8640,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df864b,
    48'h0000000df864b,
    48'h000007b034ccc,
    48'h000007b034ddc,
    48'h000007b034d71,
    48'h000007b034cb0,
    48'h000007b034c98,
    48'h000007b034c9c,
    48'h0000000df864c,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h00000423aec50,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df865a,
    48'h0000000df865a,
    48'h000007b034dfc,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h0000000df865b,
    48'h000007b034ca0,
    48'h0000040139a98,
    48'h000007b034ca0,
    48'h00000423aec50,
    48'h0000000df865c,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df865d,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df865e,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df865f,
    48'h00000423aec50,
    48'h0000000df8660,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034cba,
    48'h00000423aec50,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034dec,
    48'h000007b034de4,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb0,
    48'h000007b034d40,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb1,
    48'h000007b034d41,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ca0,
    48'h000007b034ce8,
    48'h000007b034cb2,
    48'h000007b034d42,
    48'h000007b034cba,
    48'h000007b034d4a,
    48'h000007b034cd0,
    48'h000007b034d18,
    48'h000007b034cc2,
    48'h000007b034d52,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042351e38,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df8641,
    48'h0000000df8641,
    48'h000007b034dec,
    48'h0000000df8642,
    48'h000007b034c98,
    48'h0000040139a94,
    48'h000007b034c98,
    48'h0000042351e38,
    48'h0000040138938,
    48'h0000042351e3a,
    48'h000007b034c98,
    48'h0000042351e3c,
    48'h00000400024b0,
    48'h0000040001fac,
    48'h0000000df8643,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e38,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df864d,
    48'h0000000df864d,
    48'h000007b034c9c,
    48'h0000040139a94,
    48'h000007b034c9c,
    48'h0000042351e38,
    48'h000004013893c,
    48'h0000042351e3a,
    48'h000007b034c9c,
    48'h0000042351e3c,
    48'h00000400024b0,
    48'h0000040001fac,
    48'h0000000df864e,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h00000423aec50,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df8661,
    48'h0000000df8661,
    48'h000007b034ca0,
    48'h0000040139a98,
    48'h000007b034ca0,
    48'h00000423aec50,
    48'h0000000df8662,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8663,
    48'h00000423aec50,
    48'h00000423aec54,
    48'h0000000df8664,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034dfc,
    48'h000007b034cb2,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034d94,
    48'h000004013893c,
    48'h000007b034d98,
    48'h0000040138940,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034d42,
    48'h000007b034ca0,
    48'h000007b034ce8,
    48'h000007b034cba,
    48'h000007b034d4a,
    48'h000007b034cd0,
    48'h000007b034d18,
    48'h000007b034cc2,
    48'h000007b034d52,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d30,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d42,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423aec6c,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423aec5c,
    48'h000007b034cfc,
    48'h0000040139dd8,
    48'h000007b034d98,
    48'h00000423aec60,
    48'h000007b034d00,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d42,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042351e38,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h0000042351e38,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042351e38,
    48'h0000042351e38,
    48'h0000042351e3c,
    48'h0000042351e38,
    48'h000007b034d42,
    48'h000007b034d30,
    48'h000007b034d18,
    48'h00000400015a4,
    48'h0000040138940,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h00000423aec50,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8124,
    48'h0000040136800,
    48'h00000423aec84,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423afca8,
    48'h00000423afca8,
    48'h00000423afcb4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2c8,
    48'h00000423ae400,
    48'h00000423ae400,
    48'h00000423ae40c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423afcf8,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afd08,
    48'h00000423afce8,
    48'h00000423afcec,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423afcf0,
    48'h00000423afce0,
    48'h00000423afce8,
    48'h00000423afce8,
    48'h00000423afcf0,
    48'h00000423afce0,
    48'h00000423afce8,
    48'h000004214c8a8,
    48'h00000423afd0c,
    48'h00000423afd0c,
    48'h000007b034dcc,
    48'h0000000dfcfa8,
    48'h000007b034dd4,
    48'h0000000df7c48,
    48'h000007b034dd4,
    48'h00000423afd0c,
    48'h00000423afd08,
    48'h00000423afd0c,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423afcec,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423afcf0,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df8a70,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9f10,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8a74,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000df9f14,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040136428,
    48'h000007b034a50,
    48'h000004013893c,
    48'h00000423afce0,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423afce2,
    48'h00000423afce4,
    48'h00000423afcd0,
    48'h00000423afcd0,
    48'h00000423afcd0,
    48'h00000423afcd0,
    48'h00000423afcd0,
    48'h00000423afcd4,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423afcd8,
    48'h00000423afcc8,
    48'h00000423afccc,
    48'h00000423afcd0,
    48'h00000423afcd8,
    48'h00000423afcc8,
    48'h00000423afcd4,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h00000423afcf0,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b034d58,
    48'h0000000df84d5,
    48'h000007b034dfc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354d90,
    48'h0000040138938,
    48'h0000042354d92,
    48'h000007b034c98,
    48'h0000042354d94,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h00000423afce0,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034c9c,
    48'h0000040139a84,
    48'h000007b034c9c,
    48'h00000423afce0,
    48'h0000000df84e5,
    48'h000007b034c9c,
    48'h0000040139bac,
    48'h000007b034c9c,
    48'h00000423afce0,
    48'h0000000df84e6,
    48'h000007b034c9c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034c9c,
    48'h00000423afce0,
    48'h0000000df84e7,
    48'h000007b034dfc,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h0000000df84e8,
    48'h00000423afce0,
    48'h0000000df84e9,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h0000000df84ea,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423afcec,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423afcf0,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d90,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h000007b034ce4,
    48'h000007b034d5c,
    48'h000007b034d5c,
    48'h000004013893c,
    48'h000007b034d5c,
    48'h000007b034ce4,
    48'h000007b034e94,
    48'h000007b034d5c,
    48'h000007b034dac,
    48'h000007b034e90,
    48'h000007b034d5c,
    48'h000007b034e8c,
    48'h000007b034dcc,
    48'h0000000dfb1e0,
    48'h000007b034e88,
    48'h000007b034e84,
    48'h0000040139dd4,
    48'h000007b034e90,
    48'h000007b034e8c,
    48'h000007b034e88,
    48'h000007b034e94,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce0,
    48'h00000423afce2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423afcf0,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423afcf0,
    48'h0000040022cb0,
    48'h000007b034cfc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000007b03451c,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423afcfa,
    48'h000007b034390,
    48'h000007b0344a8,
    48'h000007b034400,
    48'h000007b0344e0,
    48'h000007b034394,
    48'h000007b0344ac,
    48'h000007b034404,
    48'h000007b0344e4,
    48'h000007b034398,
    48'h000007b0344b0,
    48'h000007b034408,
    48'h000007b0344e8,
    48'h000007b03439c,
    48'h000007b0344b4,
    48'h000007b03440c,
    48'h000007b0344ec,
    48'h000007b0343a0,
    48'h000007b0344b8,
    48'h000007b034410,
    48'h000007b0344f0,
    48'h000007b0343a4,
    48'h000007b0344bc,
    48'h000007b034414,
    48'h000007b0344f4,
    48'h000007b0343a8,
    48'h000007b0344c0,
    48'h000007b034418,
    48'h000007b0344f8,
    48'h000007b0343ac,
    48'h000007b0344c4,
    48'h000007b03441c,
    48'h000007b0344fc,
    48'h000007b0343b0,
    48'h000007b0344c8,
    48'h000007b034420,
    48'h000007b034500,
    48'h000007b0343b4,
    48'h000007b0344cc,
    48'h000007b034424,
    48'h000007b034504,
    48'h000007b0343b8,
    48'h000007b0344d0,
    48'h000007b034428,
    48'h000007b034508,
    48'h000007b0343bc,
    48'h000007b0344d4,
    48'h000007b03442c,
    48'h000007b03450c,
    48'h000007b0343c0,
    48'h000007b0344d8,
    48'h000007b034430,
    48'h000007b034510,
    48'h000007b0343c4,
    48'h000007b0344dc,
    48'h000007b034434,
    48'h000007b034514,
    48'h00000423afd04,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423afd50,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afd60,
    48'h00000423afd40,
    48'h00000423afd44,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000423afd48,
    48'h00000423afd38,
    48'h00000423afd40,
    48'h00000423afd40,
    48'h00000423afd48,
    48'h00000423afd38,
    48'h00000423afd40,
    48'h000004214c8a8,
    48'h00000423afd64,
    48'h00000423afd64,
    48'h000007b034dcc,
    48'h0000000dfcfa8,
    48'h000007b034dd4,
    48'h0000000df7c48,
    48'h000007b034dd4,
    48'h00000423afd64,
    48'h00000423afd60,
    48'h00000423afd64,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423afd44,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423afd48,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df8a70,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9f10,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8a74,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000df9f14,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354d00,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040136428,
    48'h000007b034a54,
    48'h000004013893c,
    48'h00000423afd38,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423afd3a,
    48'h00000423afd3c,
    48'h00000423afd28,
    48'h00000423afd28,
    48'h00000423afd28,
    48'h00000423afd28,
    48'h00000423afd28,
    48'h00000423afd2c,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000423afd30,
    48'h00000423afd20,
    48'h00000423afd24,
    48'h00000423afd28,
    48'h00000423afd30,
    48'h00000423afd20,
    48'h00000423afd2c,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040139dd4,
    48'h00000423afd48,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354d00,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b034d58,
    48'h0000000df84d5,
    48'h000007b034dfc,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354d00,
    48'h0000040138938,
    48'h0000042354d02,
    48'h000007b034c98,
    48'h0000042354d04,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h00000423afd38,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034c9c,
    48'h0000040139a84,
    48'h000007b034c9c,
    48'h00000423afd38,
    48'h0000000df84e5,
    48'h000007b034c9c,
    48'h0000040139bac,
    48'h000007b034c9c,
    48'h00000423afd38,
    48'h0000000df84e6,
    48'h000007b034c9c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034c9c,
    48'h00000423afd38,
    48'h0000000df84e7,
    48'h000007b034dfc,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h0000000df84e8,
    48'h00000423afd38,
    48'h0000000df84e9,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h0000000df84ea,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423afd44,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423afd48,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042354d00,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h000007b034ce4,
    48'h000007b034d5c,
    48'h000007b034d5c,
    48'h000004013893c,
    48'h000007b034d5c,
    48'h000007b034ce4,
    48'h000007b034e94,
    48'h000007b034d5c,
    48'h000007b034dac,
    48'h000007b034e90,
    48'h000007b034d5c,
    48'h000007b034e8c,
    48'h000007b034dcc,
    48'h0000000dfb1e0,
    48'h000007b034e88,
    48'h000007b034e84,
    48'h0000040139dd4,
    48'h000007b034e90,
    48'h000007b034e8c,
    48'h000007b034e88,
    48'h000007b034e94,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd38,
    48'h00000423afd3a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423afd48,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423afd48,
    48'h0000040022cb0,
    48'h000007b034cfc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000007b03451c,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423afd52,
    48'h000007b034390,
    48'h000007b0344a8,
    48'h000007b034400,
    48'h000007b0344e0,
    48'h000007b034394,
    48'h000007b0344ac,
    48'h000007b034404,
    48'h000007b0344e4,
    48'h000007b034398,
    48'h000007b0344b0,
    48'h000007b034408,
    48'h000007b0344e8,
    48'h000007b03439c,
    48'h000007b0344b4,
    48'h000007b03440c,
    48'h000007b0344ec,
    48'h000007b0343a0,
    48'h000007b0344b8,
    48'h000007b034410,
    48'h000007b0344f0,
    48'h000007b0343a4,
    48'h000007b0344bc,
    48'h000007b034414,
    48'h000007b0344f4,
    48'h000007b0343a8,
    48'h000007b0344c0,
    48'h000007b034418,
    48'h000007b0344f8,
    48'h000007b0343ac,
    48'h000007b0344c4,
    48'h000007b03441c,
    48'h000007b0344fc,
    48'h000007b0343b0,
    48'h000007b0344c8,
    48'h000007b034420,
    48'h000007b034500,
    48'h000007b0343b4,
    48'h000007b0344cc,
    48'h000007b034424,
    48'h000007b034504,
    48'h000007b0343b8,
    48'h000007b0344d0,
    48'h000007b034428,
    48'h000007b034508,
    48'h000007b0343bc,
    48'h000007b0344d4,
    48'h000007b03442c,
    48'h000007b03450c,
    48'h000007b0343c0,
    48'h000007b0344d8,
    48'h000007b034430,
    48'h000007b034510,
    48'h000007b0343c4,
    48'h000007b0344dc,
    48'h000007b034434,
    48'h000007b034514,
    48'h00000423afd5c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423afda8,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afdb8,
    48'h00000423afd80,
    48'h00000423afd84,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423afd88,
    48'h00000423afd70,
    48'h00000423afd80,
    48'h00000423afd80,
    48'h00000423afd88,
    48'h00000423afd70,
    48'h00000423afd80,
    48'h000004214c8a8,
    48'h00000423afdbc,
    48'h00000423afdbc,
    48'h000007b034dcc,
    48'h0000000dfd064,
    48'h000007b034dd4,
    48'h0000000df7d04,
    48'h000007b034dd4,
    48'h00000423afdbc,
    48'h00000423afdb8,
    48'h00000423afdbc,
    48'h00000400026f0,
    48'h0000040139dd0,
    48'h00000423afd84,
    48'h0000040138938,
    48'h00000423afd88,
    48'h0000040139dd4,
    48'h00000423afd74,
    48'h000004013893c,
    48'h00000423afd88,
    48'h0000040139dd8,
    48'h00000423afd78,
    48'h0000040138940,
    48'h000007b034dcc,
    48'h0000000df8e1c,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000dfa2bc,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8e20,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000dfa2c0,
    48'h000007b034dac,
    48'h000007b034dcc,
    48'h0000000df8e24,
    48'h000007b034c58,
    48'h000007b034c70,
    48'h0000000dfa2c4,
    48'h000007b034db0,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df863c,
    48'h0000000df863d,
    48'h0000000df863e,
    48'h0000000df863f,
    48'h0000000df8640,
    48'h0000000df8641,
    48'h0000000df8642,
    48'h0000000df8643,
    48'h0000000df8644,
    48'h0000000df8645,
    48'h0000000df8646,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df8648,
    48'h0000000df8649,
    48'h0000040138938,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034d71,
    48'h0000040138938,
    48'h0000040138940,
    48'h0000042354e20,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h000007b034d72,
    48'h0000000df864a,
    48'h0000000df864b,
    48'h0000040138938,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034d71,
    48'h0000040138938,
    48'h0000040138940,
    48'h0000042354e20,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h000007b034d72,
    48'h0000000df864c,
    48'h0000000df864d,
    48'h0000000df864e,
    48'h0000000df864f,
    48'h0000000df8650,
    48'h0000000df8651,
    48'h0000000df8652,
    48'h0000040138940,
    48'h000007b034d98,
    48'h000007b034c70,
    48'h0000000df8654,
    48'h0000000df8655,
    48'h0000000df8656,
    48'h0000000df8657,
    48'h0000000df8658,
    48'h0000000df8659,
    48'h0000000df865a,
    48'h0000000df865b,
    48'h0000000df865c,
    48'h0000000df865d,
    48'h0000000df865e,
    48'h0000000df865f,
    48'h0000000df8660,
    48'h0000000df8661,
    48'h0000000df8662,
    48'h0000000df8663,
    48'h0000000df8664,
    48'h0000000df8665,
    48'h0000000df8666,
    48'h0000040138938,
    48'h0000042354e20,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df863c,
    48'h0000040138938,
    48'h0000042354e24,
    48'h00000401367d0,
    48'h000007b0345b4,
    48'h0000040136428,
    48'h000007b034a34,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df8648,
    48'h000004013893c,
    48'h0000042354e24,
    48'h00000401367d0,
    48'h000007b0345b4,
    48'h0000040136428,
    48'h000007b034a34,
    48'h0000040138940,
    48'h0000042351e00,
    48'h000007b034d60,
    48'h000007b034c88,
    48'h000007b034c70,
    48'h0000000df8654,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354e20,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df863c,
    48'h0000000df863c,
    48'h000007b034d58,
    48'h0000000df863d,
    48'h000007b034dfc,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000000df863e,
    48'h000007b034c68,
    48'h000007b034cc0,
    48'h000007b034cb8,
    48'h000007b034de4,
    48'h0000042354e20,
    48'h000007b034c98,
    48'h000007b034cc8,
    48'h000007b034de4,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df8648,
    48'h0000000df8648,
    48'h0000000df8649,
    48'h000007b034ccc,
    48'h000007b034ddc,
    48'h000007b034d71,
    48'h000007b034cb0,
    48'h000007b034c98,
    48'h000007b034c9c,
    48'h0000000df864a,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034cb9,
    48'h0000042354e20,
    48'h000007b034c9c,
    48'h000007b034ccc,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h0000042351e00,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df8654,
    48'h0000000df8654,
    48'h000007b034ca0,
    48'h0000040139a84,
    48'h000007b034ca0,
    48'h0000042351e00,
    48'h0000000df8655,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df8656,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df8657,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df8658,
    48'h0000042351e00,
    48'h0000000df8659,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034dfc,
    48'h000007b034cb2,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034dec,
    48'h000007b034de4,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354e20,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df863f,
    48'h0000000df863f,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354e20,
    48'h0000040138938,
    48'h0000042354e22,
    48'h000007b034c98,
    48'h0000042354e24,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df8640,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df864b,
    48'h0000000df864b,
    48'h000007b034ccc,
    48'h000007b034ddc,
    48'h000007b034d71,
    48'h000007b034cb0,
    48'h000007b034c98,
    48'h000007b034c9c,
    48'h0000000df864c,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c70,
    48'h0000040138940,
    48'h0000042351e00,
    48'h000007b034ca0,
    48'h000007b034cb2,
    48'h000007b034cba,
    48'h000007b034cc2,
    48'h000007b034cd0,
    48'h0000000df865a,
    48'h0000000df865a,
    48'h000007b034dfc,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000000df865b,
    48'h000007b034ca0,
    48'h0000040139a98,
    48'h000007b034ca0,
    48'h0000042351e00,
    48'h0000000df865c,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df865d,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df865e,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df865f,
    48'h0000042351e00,
    48'h0000000df8660,
    48'h000007b034c70,
    48'h000007b034ca0,
    48'h000007b034cc2,
    48'h000007b034dfc,
    48'h000007b034cb2,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034cc2,
    48'h000007b034d94,
    48'h000004013893c,
    48'h000007b034d98,
    48'h0000040138940,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034d42,
    48'h000007b034ca0,
    48'h000007b034ce8,
    48'h000007b034cba,
    48'h000007b034d4a,
    48'h000007b034cd0,
    48'h000007b034d18,
    48'h000007b034cc2,
    48'h000007b034d52,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d30,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d42,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423afd84,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423afd74,
    48'h000007b034cfc,
    48'h0000040139dd8,
    48'h000007b034d98,
    48'h00000423afd78,
    48'h000007b034d00,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d42,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e20,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h000007b034d42,
    48'h000007b034d30,
    48'h000007b034d18,
    48'h00000400015a4,
    48'h0000040138940,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8124,
    48'h0000040136800,
    48'h00000423afdb4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423ae428,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423ae438,
    48'h00000423ae418,
    48'h00000423ae41c,
    48'h0000042351df0,
    48'h00000423ae418,
    48'h00000423ae418,
    48'h00000423ae420,
    48'h0000042354d90,
    48'h00000423ae418,
    48'h000004214c8a8,
    48'h00000423ae43c,
    48'h00000423ae43c,
    48'h000007b034dcc,
    48'h0000000dfcf34,
    48'h000007b034dd4,
    48'h0000000df7bd4,
    48'h000007b034dd4,
    48'h00000423ae43c,
    48'h00000423ae438,
    48'h00000423ae43c,
    48'h00000400025c0,
    48'h0000040139dd0,
    48'h00000423ae420,
    48'h0000040138938,
    48'h000007b034dcc,
    48'h0000000df882c,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9ccc,
    48'h000007b034da8,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df8420,
    48'h0000000df8421,
    48'h0000000df8422,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df8420,
    48'h0000040138938,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040136428,
    48'h000007b034a50,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df8420,
    48'h0000000df8420,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354d90,
    48'h0000040138938,
    48'h0000042354d92,
    48'h000007b034c98,
    48'h0000042354d94,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df8421,
    48'h000007b034dfc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000000df8422,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034cc0,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d40,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423ae420,
    48'h000007b034cf8,
    48'h000007b034d40,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d90,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df7ff4,
    48'h0000040136800,
    48'h00000423ae434,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423ae498,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423ae4a8,
    48'h00000423ae488,
    48'h00000423ae48c,
    48'h0000042351de8,
    48'h00000423ae488,
    48'h00000423ae488,
    48'h00000423ae490,
    48'h00000423ae478,
    48'h00000423ae488,
    48'h000004214c8a8,
    48'h00000423ae4ac,
    48'h00000423ae4ac,
    48'h000007b034dcc,
    48'h0000000dfd28c,
    48'h000007b034dd4,
    48'h0000000df7f2c,
    48'h000007b034dd4,
    48'h0000040136800,
    48'h00000423ae4a4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423afe90,
    48'h00000423afe90,
    48'h00000423afe9c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2cc,
    48'h00000423b0050,
    48'h00000423b0050,
    48'h00000423b005c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2d0,
    48'h00000423afeb8,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afec8,
    48'h00000423afea8,
    48'h00000423afeac,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h00000423afeb0,
    48'h0000042351e00,
    48'h00000423afea8,
    48'h00000423afea8,
    48'h00000423afeb0,
    48'h0000042351e00,
    48'h00000423afea8,
    48'h000004214c8a8,
    48'h00000423afecc,
    48'h00000423afecc,
    48'h000007b034dcc,
    48'h0000000dfcfa8,
    48'h000007b034dd4,
    48'h0000000df7c48,
    48'h000007b034dd4,
    48'h00000423afecc,
    48'h00000423afec8,
    48'h00000423afecc,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423afeac,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423afeb0,
    48'h000004013893c,
    48'h000007b034dcc,
    48'h0000000df8a70,
    48'h000007b034c50,
    48'h000007b034c68,
    48'h0000000df9f10,
    48'h000007b034da8,
    48'h000007b034dcc,
    48'h0000000df8a74,
    48'h000007b034c54,
    48'h000007b034c6c,
    48'h0000000df9f14,
    48'h000007b034dac,
    48'h0000040138938,
    48'h000007b034d90,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b034d94,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354c70,
    48'h000007b034d58,
    48'h000007b034c80,
    48'h000007b034c68,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354c74,
    48'h00000401367d0,
    48'h000007b0345a8,
    48'h0000040136428,
    48'h000007b034a28,
    48'h000004013893c,
    48'h0000042351e00,
    48'h000007b034d5c,
    48'h000007b034c84,
    48'h000007b034c6c,
    48'h0000000df84e4,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354c70,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b034d58,
    48'h0000000df84d5,
    48'h000007b034dfc,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h000007b034c98,
    48'h0000040139a98,
    48'h000007b034c98,
    48'h0000042354c70,
    48'h0000040138938,
    48'h0000042354c72,
    48'h000007b034c98,
    48'h0000042354c74,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e00,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034c9c,
    48'h0000040139a84,
    48'h000007b034c9c,
    48'h0000042351e00,
    48'h0000000df84e5,
    48'h000007b034c9c,
    48'h0000040139bac,
    48'h000007b034c9c,
    48'h0000042351e00,
    48'h0000000df84e6,
    48'h000007b034c9c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034c9c,
    48'h0000042351e00,
    48'h0000000df84e7,
    48'h000007b034dfc,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000000df84e8,
    48'h0000042351e00,
    48'h0000042351e04,
    48'h0000000df84e9,
    48'h0000042351e00,
    48'h0000000df84ea,
    48'h000007b034c6c,
    48'h000007b034c9c,
    48'h000007b034cc1,
    48'h000007b034cb9,
    48'h0000042351e00,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034dec,
    48'h000007b034de4,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb0,
    48'h000007b034d40,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb1,
    48'h000007b034d41,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034dd4,
    48'h000007b034de4,
    48'h000007b034dec,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c68,
    48'h0000040138938,
    48'h0000042354c70,
    48'h000007b034c98,
    48'h000007b034cb0,
    48'h000007b034cb8,
    48'h000007b034cc0,
    48'h000007b034cc8,
    48'h0000000df84d7,
    48'h0000000df84d7,
    48'h000007b034c98,
    48'h0000040139a84,
    48'h000007b034c98,
    48'h0000042354c70,
    48'h0000040138938,
    48'h0000042354c72,
    48'h000007b034c98,
    48'h0000042354c74,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df84d8,
    48'h000007b034c98,
    48'h0000040139bac,
    48'h000007b034c98,
    48'h0000042354c70,
    48'h0000040138938,
    48'h0000042354c72,
    48'h000007b034c98,
    48'h0000042354c74,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d9,
    48'h000007b034c68,
    48'h000007b034c98,
    48'h000007b034cc0,
    48'h000007b034dfc,
    48'h000007b034cb0,
    48'h000007b034dfc,
    48'h000007b034df4,
    48'h000007b034c6c,
    48'h000004013893c,
    48'h0000042351e00,
    48'h000007b034c9c,
    48'h000007b034cb1,
    48'h000007b034cb9,
    48'h000007b034cc1,
    48'h000007b034ccc,
    48'h0000000df84eb,
    48'h0000000df84eb,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000000df84ec,
    48'h000007b034c6c,
    48'h000007b034cc1,
    48'h000007b034dfc,
    48'h000007b034cb1,
    48'h000007b034cc0,
    48'h000007b034cc1,
    48'h000007b034d40,
    48'h000007b034c98,
    48'h000007b034ce0,
    48'h000007b034cb8,
    48'h000007b034d48,
    48'h000007b034cc8,
    48'h000007b034d10,
    48'h000007b034cc0,
    48'h000007b034d50,
    48'h000007b034d41,
    48'h000007b034c9c,
    48'h000007b034ce4,
    48'h000007b034cb9,
    48'h000007b034d49,
    48'h000007b034ccc,
    48'h000007b034d14,
    48'h000007b034cc1,
    48'h000007b034d51,
    48'h000007b034ddc,
    48'h000007b034d28,
    48'h000007b034d2c,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h0000040139dd0,
    48'h000007b034d90,
    48'h00000423afeac,
    48'h000007b034cf8,
    48'h0000040139dd4,
    48'h000007b034d94,
    48'h00000423afeb0,
    48'h000007b034cfc,
    48'h000007b034d40,
    48'h000007b034d41,
    48'h000007b034d40,
    48'h000007b034d28,
    48'h000007b034d10,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h0000042354c70,
    48'h000007b034d41,
    48'h000007b034d2c,
    48'h000007b034d14,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000042351e00,
    48'h0000040136800,
    48'h000007b034dcc,
    48'h0000000df8068,
    48'h0000040136800,
    48'h00000423afec4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2d0,
    48'h00000423afee0,
    48'h000007b0344a8,
    48'h000007b0344e0,
    48'h000007b0344ac,
    48'h000007b0344e4,
    48'h000007b0344b0,
    48'h000007b0344e8,
    48'h000007b0344b4,
    48'h000007b0344ec,
    48'h000007b0344b8,
    48'h000007b0344f0,
    48'h000007b0344bc,
    48'h000007b0344f4,
    48'h000007b0344c0,
    48'h000007b0344f8,
    48'h000007b0344c4,
    48'h000007b0344fc,
    48'h000007b0344c8,
    48'h000007b034500,
    48'h000007b0344cc,
    48'h000007b034504,
    48'h000007b0344d0,
    48'h000007b034508,
    48'h000007b0344d4,
    48'h000007b03450c,
    48'h000007b0344d8,
    48'h000007b034510,
    48'h000007b0344dc,
    48'h000007b034514,
    48'h0000040023c88,
    48'h000007b034c14,
    48'h000007b034dc4,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034c14,
    48'h0000040022e78,
    48'h00000423afef0,
    48'h00000423afed8,
    48'h0000040136800,
    48'h00000423afeec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2d0,
    48'h00000423aff58,
    48'h00000423aff58,
    48'h00000423aff64,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af2d0,
    48'h0000042354c78,
    48'h0000042354c78,
    48'h0000042354c84,
    48'h000007b0343c8,
    48'h000007b0343cc,
    48'h000007b0343d0,
    48'h000007b0343d4,
    48'h000007b0343d8,
    48'h000007b0343dc,
    48'h000007b0343e0,
    48'h000007b0343e4,
    48'h000007b0343e8,
    48'h000007b0343ec,
    48'h000007b0343f0,
    48'h000007b0343f4,
    48'h000007b0343f8,
    48'h000007b0343fc,
    48'h0000040023890,
    48'h000007b034390,
    48'h000007b034400,
    48'h000007b034438,
    48'h000007b034394,
    48'h000007b034404,
    48'h000007b03443c,
    48'h000007b034398,
    48'h000007b034408,
    48'h000007b034440,
    48'h000007b03439c,
    48'h000007b03440c,
    48'h000007b034444,
    48'h000007b0343a0,
    48'h000007b034410,
    48'h000007b034448,
    48'h000007b0343a4,
    48'h000007b034524,
    48'h0000040023890,
    48'h000007b034400,
    48'h000007b034390,
    48'h000007b034438,
    48'h000007b034404,
    48'h000007b034394,
    48'h000007b03443c,
    48'h000007b034408,
    48'h000007b034398,
    48'h000007b034440,
    48'h000007b03440c,
    48'h000007b03439c,
    48'h000007b034444,
    48'h000007b034410,
    48'h000007b0343a0,
    48'h000007b034448,
    48'h000007b034414,
    48'h000007b0343a4,
    48'h0000040023b70,
    48'h0000040002490,
    48'h000007b034c14,
    48'h000007b034c10,
    48'h0000040023b70,
    48'h000007b034c10,
    48'h0000040023b70,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040023892,
    48'h0000040023a5a,
    48'h0000040023aca,
    48'h000007b0343a4,
    48'h000007b0343a4,
    48'h0000040139780,
    48'h0000040139780,
    48'h000007b0343a8,
    48'h000007b0343a8,
    48'h0000040139784,
    48'h0000040139784,
    48'h000007b0343ac,
    48'h000007b0343ac,
    48'h0000040139788,
    48'h0000040139788,
    48'h000007b0343b0,
    48'h000007b0343b0,
    48'h000004013978c,
    48'h000004013978c,
    48'h000007b0343b8,
    48'h000007b0343b8,
    48'h0000040139790,
    48'h0000040139790,
    48'h000007b0343bc,
    48'h000007b0343bc,
    48'h0000040139794,
    48'h0000040139794,
    48'h000007b0343c0,
    48'h000007b0343c0,
    48'h0000040139798,
    48'h0000040139798,
    48'h000007b0343c4,
    48'h000007b0343c4,
    48'h000004013979c,
    48'h000007b03444c,
    48'h000007b034c14,
    48'h0000040023890,
    48'h0000040023b38,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc0,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc2,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc4,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc6,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbc8,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbca,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbcc,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbce,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd0,
    48'h0000040139068,
    48'h0000042352bd0,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd2,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd4,
    48'h0000040139068,
    48'h0000042352bd8,
    48'h00000423ace3a,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd6,
    48'h0000040139068,
    48'h0000042352bdc,
    48'h00000423aceca,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbd8,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbda,
    48'h0000040139068,
    48'h0000042352be4,
    48'h00000423ad2ca,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbdc,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbde,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe0,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe2,
    48'h0000040139068,
    48'h0000042352bf4,
    48'h00000423adaea,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe4,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe6,
    48'h0000040139068,
    48'h0000042352bfc,
    48'h00000423ae05a,
    48'h0000040001fac,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbe8,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbea,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbec,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbee,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbf0,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbf2,
    48'h000004214c578,
    48'h0000040138950,
    48'h00000423afbf4,
    48'h000004214c578,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040023890,
    48'h0000040138b29,
    48'h000007b0343a4,
    48'h000007b03444c,
    48'h000007b034418,
    48'h000007b0343a8,
    48'h000007b034450,
    48'h000007b03441c,
    48'h000007b0343ac,
    48'h000007b034454,
    48'h000007b034420,
    48'h000007b0343b0,
    48'h000007b034458,
    48'h000007b034424,
    48'h000007b0343b4,
    48'h000007b03445c,
    48'h000007b034428,
    48'h000007b0343b8,
    48'h000007b034460,
    48'h000007b03442c,
    48'h000007b0343bc,
    48'h000007b034464,
    48'h000007b034430,
    48'h000007b0343c0,
    48'h000007b034468,
    48'h000007b034434,
    48'h000007b0343c4,
    48'h000007b03446c,
    48'h000004213c268,
    48'h0000040139038,
    48'h000007b03451c,
    48'h000004214c578,
    48'h0000040023760,
    48'h000004214c578,
    48'h0000040023768,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h0000042354b84,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354b78,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354b7a,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h0000042354b88,
    48'h0000042354b68,
    48'h0000042354b6c,
    48'h0000042354b60,
    48'h0000042354b64,
    48'h0000042354b70,
    48'h0000042354af8,
    48'h0000042354b68,
    48'h0000042354b68,
    48'h0000042354b70,
    48'h0000042354af8,
    48'h0000042354b68,
    48'h000004214c8a8,
    48'h0000042354b8c,
    48'h0000042354b8c,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h0000042354b8c,
    48'h0000042354b88,
    48'h0000042354b8c,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h0000042354b6c,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042354b70,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354b60,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354b64,
    48'h00000401367d0,
    48'h000007b0345c0,
    48'h0000040136428,
    48'h000007b034a40,
    48'h000004013893c,
    48'h0000042354af8,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h0000042354afa,
    48'h0000042354afc,
    48'h0000042354ae8,
    48'h0000042354ae8,
    48'h0000042354ae8,
    48'h0000042354ae8,
    48'h0000042354ae8,
    48'h0000042354aec,
    48'h0000042351e40,
    48'h0000042351e44,
    48'h0000042354af0,
    48'h0000042354ae0,
    48'h0000042354ae4,
    48'h0000042354ae8,
    48'h0000042354af0,
    48'h0000042354ae0,
    48'h0000042354aec,
    48'h0000042351e40,
    48'h0000042351e44,
    48'h00000401367d0,
    48'h000007b0345e0,
    48'h0000040139dd4,
    48'h0000042354b70,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042354b60,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042354b60,
    48'h0000042354b64,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042354b60,
    48'h0000040138938,
    48'h0000042354b62,
    48'h000007b034f58,
    48'h0000042354b64,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042354af8,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042354af8,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042354af8,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042354af8,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000000df84e8,
    48'h0000042354af8,
    48'h0000000df84e9,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h0000042354b6c,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042354b70,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354b60,
    48'h0000042354b60,
    48'h0000042354b64,
    48'h0000042354b60,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354af8,
    48'h0000042354afa,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042354b70,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042354b70,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034ba8,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000042354b88,
    48'h0000042354b68,
    48'h0000042354b6c,
    48'h0000042354b60,
    48'h0000042354b60,
    48'h0000042354b60,
    48'h0000042354b64,
    48'h0000042354b62,
    48'h0000040001fac,
    48'h0000040023a64,
    48'h0000040023768,
    48'h000007b034e2e,
    48'h0000040023760,
    48'h000007b034cc0,
    48'h0000042354b94,
    48'h0000042354b9a,
    48'h0000042354ba0,
    48'h0000042354b78,
    48'h0000042354b78,
    48'h000004213c310,
    48'h0000042354c4c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354c40,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354c42,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h0000042354c50,
    48'h0000042354c30,
    48'h0000042354c34,
    48'h0000042354c28,
    48'h0000042354c2c,
    48'h0000042354c38,
    48'h0000042354bc0,
    48'h0000042354c30,
    48'h0000042354c30,
    48'h0000042354c38,
    48'h0000042354bc0,
    48'h0000042354c30,
    48'h000004214c8a8,
    48'h0000042354c54,
    48'h0000042354c54,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h0000042354c54,
    48'h0000042354c50,
    48'h0000042354c54,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h0000042354c34,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042354c38,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354c28,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354c2c,
    48'h00000401367d0,
    48'h000007b0345bc,
    48'h0000040136428,
    48'h000007b034a3c,
    48'h000004013893c,
    48'h0000042354bc0,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h0000042354bc2,
    48'h0000042354bc4,
    48'h0000042354bb0,
    48'h0000042354bb0,
    48'h0000042354bb0,
    48'h0000042354bb0,
    48'h0000042354bb0,
    48'h0000042354bb4,
    48'h0000042351e40,
    48'h0000042351e44,
    48'h0000042354bb8,
    48'h0000042354ba8,
    48'h0000042354bac,
    48'h0000042354bb0,
    48'h0000042354bb8,
    48'h0000042354ba8,
    48'h0000042354bb4,
    48'h0000042351e40,
    48'h0000042351e44,
    48'h00000401367d0,
    48'h000007b0345e0,
    48'h0000040139dd4,
    48'h0000042354c38,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042354c28,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042354c28,
    48'h0000042354c2c,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042354c28,
    48'h0000040138938,
    48'h0000042354c2a,
    48'h000007b034f58,
    48'h0000042354c2c,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042354bc0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042354bc0,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042354bc0,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042354bc0,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000000df84e8,
    48'h0000042354bc0,
    48'h0000000df84e9,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h0000042354c34,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042354c38,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354c28,
    48'h0000042354c28,
    48'h0000042354c2c,
    48'h0000042354c28,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc0,
    48'h0000042354bc2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042354c38,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042354c38,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034ba8,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000042354c50,
    48'h0000042354c30,
    48'h0000042354c34,
    48'h0000042354c28,
    48'h0000042354c28,
    48'h0000042354c28,
    48'h0000042354c2c,
    48'h0000042354c2a,
    48'h0000040001fac,
    48'h0000040023a62,
    48'h0000040023768,
    48'h000007b034e2d,
    48'h0000040023760,
    48'h000007b034cbc,
    48'h0000042354c5c,
    48'h0000042354c62,
    48'h0000042354c68,
    48'h0000042354c40,
    48'h0000042354c40,
    48'h000004213c310,
    48'h0000042354c9c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354c90,
    48'h0000042354c90,
    48'h0000042354c90,
    48'h0000042354c90,
    48'h000004213c310,
    48'h0000042354d24,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354d18,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354d1a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042354d28,
    48'h0000042354d08,
    48'h0000042354d0c,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042354d02,
    48'h0000040001fac,
    48'h0000040023a6e,
    48'h0000040023768,
    48'h000007b034e33,
    48'h0000040023760,
    48'h000007b034cd4,
    48'h0000042354d34,
    48'h0000042354d18,
    48'h0000042354d18,
    48'h000004213c310,
    48'h0000042354db4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354da8,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354daa,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042354db8,
    48'h0000042354d98,
    48'h0000042354d9c,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d92,
    48'h0000040001fac,
    48'h0000040023a6c,
    48'h0000040023768,
    48'h000007b034e32,
    48'h0000040023760,
    48'h000007b034cd0,
    48'h0000042354dc4,
    48'h0000042354da8,
    48'h0000042354da8,
    48'h000004213c310,
    48'h0000042354ebc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354eb0,
    48'h0000042354eb0,
    48'h0000042354eb0,
    48'h0000042354eb0,
    48'h000004213c310,
    48'h0000042354eec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354ee0,
    48'h0000042354ee0,
    48'h0000042354ee0,
    48'h0000042354ee0,
    48'h000004213c310,
    48'h0000042354f1c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354f10,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354f12,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042354f20,
    48'h0000042354f00,
    48'h0000042354f04,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h0000040023a5e,
    48'h0000040023768,
    48'h000007b034e2b,
    48'h0000040023760,
    48'h000007b034cb4,
    48'h0000042354f2c,
    48'h0000042354f10,
    48'h0000042354f10,
    48'h000004213c310,
    48'h00000423b032c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h00000423b0320,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423b0322,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423b0330,
    48'h00000423b0310,
    48'h00000423b0314,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h00000423b033c,
    48'h00000423b0320,
    48'h00000423b0320,
    48'h000004213c310,
    48'h00000423b03a4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h00000423b0398,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423b039a,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423b03a8,
    48'h00000423b0358,
    48'h00000423b035c,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h00000423b03b4,
    48'h00000423b0398,
    48'h00000423b0398,
    48'h000004213c310,
    48'h0000042354f6c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042354f60,
    48'h0000042354f60,
    48'h0000042354f60,
    48'h0000042354f60,
    48'h000004213c310,
    48'h00000423557a4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af25c,
    48'h0000042355798,
    48'h0000042355798,
    48'h0000042355798,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042355798,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h0000042355054,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af260,
    48'h0000042355048,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235504a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042355064,
    48'h0000042355048,
    48'h0000042355048,
    48'h000004213c310,
    48'h00000423550c4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af260,
    48'h00000423550b8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423550ba,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423550c8,
    48'h00000423550a8,
    48'h00000423550ac,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h00000423550d4,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h000004213c310,
    48'h00000423550ec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af260,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h000004213c310,
    48'h000004235515c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af260,
    48'h0000042355150,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355152,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h000004235513c,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355140,
    48'h0000042355140,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355140,
    48'h000004214c8a8,
    48'h0000042355164,
    48'h0000042355164,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h0000042355164,
    48'h0000042355160,
    48'h0000042355164,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h0000042355144,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042355148,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042355138,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h000004235513c,
    48'h00000401367d0,
    48'h000007b0345c8,
    48'h0000040136428,
    48'h000007b034a48,
    48'h000004013893c,
    48'h0000042355130,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h0000042355132,
    48'h0000042355134,
    48'h0000042355120,
    48'h0000042355120,
    48'h0000042355120,
    48'h0000042355120,
    48'h0000042355120,
    48'h0000042355124,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042355128,
    48'h0000042355118,
    48'h000004235511c,
    48'h0000042355120,
    48'h0000042355128,
    48'h0000042355118,
    48'h0000042355124,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040139dd4,
    48'h0000042355148,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355138,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042355138,
    48'h000004235513c,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042355138,
    48'h0000040138938,
    48'h000004235513a,
    48'h000007b034f58,
    48'h000004235513c,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042355130,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042355130,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042355130,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042355130,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000000df84e8,
    48'h0000042355130,
    48'h0000000df84e9,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h0000042355144,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042355148,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042355138,
    48'h0000042355138,
    48'h000004235513c,
    48'h0000042355138,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355130,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355132,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042355148,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042355148,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034baa,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c780,
    48'h0000040139978,
    48'h000004214c490,
    48'h0000042355130,
    48'h0000040138f40,
    48'h0000042355130,
    48'h000004214c490,
    48'h0000040139978,
    48'h000004214c698,
    48'h0000042355130,
    48'h0000042355130,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c490,
    48'h0000040139540,
    48'h000007b035194,
    48'h0000042355130,
    48'h0000042355130,
    48'h0000042355134,
    48'h0000042355130,
    48'h0000042355120,
    48'h00000400015bc,
    48'h0000042355158,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e8,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h00000423550c0,
    48'h0000042355048,
    48'h0000042355048,
    48'h000007b035154,
    48'h000004235504c,
    48'h000004213a120,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042355040,
    48'h0000042354d90,
    48'h000004235503c,
    48'h0000042355130,
    48'h0000042351df0,
    48'h0000042355050,
    48'h0000042355798,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000007b034fb8,
    48'h0000040139978,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h0000042355138,
    48'h0000042355138,
    48'h000004235513c,
    48'h000004235513a,
    48'h0000040001fac,
    48'h0000040023a68,
    48'h0000040023768,
    48'h000007b034e30,
    48'h0000040023760,
    48'h000007b034cc8,
    48'h000004235516c,
    48'h0000042355150,
    48'h0000042355150,
    48'h000004213c310,
    48'h00000423551ec,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af264,
    48'h00000423551e0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423551e2,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423551f0,
    48'h00000423551d0,
    48'h00000423551d4,
    48'h0000042351df0,
    48'h00000423551d0,
    48'h00000423551d0,
    48'h00000423551d8,
    48'h00000423551c0,
    48'h00000423551d0,
    48'h000004214c8a8,
    48'h00000423551f4,
    48'h00000423551f4,
    48'h000007b03508c,
    48'h0000000dfcf58,
    48'h000007b035094,
    48'h0000000df7bf8,
    48'h000007b035094,
    48'h00000423551f4,
    48'h00000423551f0,
    48'h00000423551f4,
    48'h00000400025e4,
    48'h00000423551d8,
    48'h0000040139dd0,
    48'h00000423551c4,
    48'h0000040138938,
    48'h00000423551d8,
    48'h0000040139dd4,
    48'h00000423551c8,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df88e0,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9d80,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df88e4,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9d84,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df8444,
    48'h0000000df8445,
    48'h0000000df8446,
    48'h0000000df8447,
    48'h0000000df8448,
    48'h0000000df8449,
    48'h0000000df844a,
    48'h0000000df844b,
    48'h0000000df844c,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df8450,
    48'h0000000df8451,
    48'h0000000df8452,
    48'h0000000df8453,
    48'h0000000df8454,
    48'h0000000df8455,
    48'h0000000df8456,
    48'h0000000df8457,
    48'h0000000df8458,
    48'h0000040138938,
    48'h0000042355190,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df8444,
    48'h0000040138938,
    48'h0000040139dd0,
    48'h0000042355192,
    48'h0000042355194,
    48'h0000042355180,
    48'h0000042355180,
    48'h0000042355180,
    48'h0000042355180,
    48'h0000042355180,
    48'h0000042355184,
    48'h0000042355138,
    48'h000004235513c,
    48'h0000042355188,
    48'h0000042355178,
    48'h000004235517c,
    48'h0000042355180,
    48'h0000042355188,
    48'h0000042355178,
    48'h0000042355184,
    48'h0000042355138,
    48'h000004235513c,
    48'h00000401367d0,
    48'h000007b0345c8,
    48'h0000040139dd0,
    48'h00000423551c4,
    48'h0000040138938,
    48'h000007b035050,
    48'h000004013893c,
    48'h00000423551b8,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df8450,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423551ba,
    48'h00000423551bc,
    48'h00000423551a8,
    48'h00000423551a8,
    48'h00000423551a8,
    48'h00000423551a8,
    48'h00000423551a8,
    48'h00000423551ac,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423551b0,
    48'h00000423551a0,
    48'h00000423551a4,
    48'h00000423551a8,
    48'h00000423551b0,
    48'h00000423551a0,
    48'h00000423551ac,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h00000423551c8,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355190,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df8444,
    48'h0000000df8444,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042355190,
    48'h0000000df8445,
    48'h0000042355190,
    48'h0000000df8446,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000000df8447,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h0000042355190,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423551b8,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8450,
    48'h0000000df8450,
    48'h000007b0350bc,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h0000000df8451,
    48'h000007b034f5c,
    48'h0000040139a98,
    48'h000007b034f5c,
    48'h00000423551b8,
    48'h0000000df8452,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355190,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df8448,
    48'h0000000df8448,
    48'h000007b0350bc,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000000df8449,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042355190,
    48'h0000000df844a,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423551b8,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8453,
    48'h0000000df8453,
    48'h00000423551b8,
    48'h0000000df8454,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h0000000df8455,
    48'h000007b034f5c,
    48'h0000040139a98,
    48'h000007b034f5c,
    48'h00000423551b8,
    48'h0000000df8456,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423551b8,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355190,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df844b,
    48'h0000000df844b,
    48'h0000042355190,
    48'h000007b034f40,
    48'h0000042355194,
    48'h0000042355180,
    48'h0000000df844c,
    48'h000007b034f28,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h000007b0350a4,
    48'h0000042355190,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423551b8,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8457,
    48'h0000000df8457,
    48'h00000423551b8,
    48'h000007b034f44,
    48'h00000423551bc,
    48'h00000423551a8,
    48'h0000000df8458,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h000007b0350a4,
    48'h00000423551b8,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b034fd0,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423551c4,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423551c8,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h0000040138938,
    48'h0000042355190,
    48'h0000042355190,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fd0,
    48'h000007b034fe8,
    48'h000007b035008,
    48'h000007b034fe8,
    48'h000007b035018,
    48'h0000040138938,
    48'h000007b035018,
    48'h000007b034fa0,
    48'h000007b035154,
    48'h000007b035018,
    48'h000007b035068,
    48'h000007b035150,
    48'h000007b035018,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb17b,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd0,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355192,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423551c4,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423551c4,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fb8,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb17c,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551ba,
    48'h0000040136800,
    48'h0000040139540,
    48'h000004214c780,
    48'h000004214c490,
    48'h0000042355190,
    48'h0000042355190,
    48'h00000423551b8,
    48'h0000042355192,
    48'h00000423551ba,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h0000042355194,
    48'h00000423551bc,
    48'h0000042355180,
    48'h00000423551a8,
    48'h0000042355182,
    48'h00000423551aa,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h0000042355188,
    48'h00000423551b0,
    48'h0000042355178,
    48'h00000423551a0,
    48'h000004235517a,
    48'h00000423551a2,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h000004235517c,
    48'h00000423551a4,
    48'h00000003840fc,
    48'h0000042355184,
    48'h00000423551ac,
    48'h0000042355138,
    48'h0000042354d90,
    48'h000004235513a,
    48'h0000042354d92,
    48'h000004235513c,
    48'h0000042354d94,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040139540,
    48'h000004214c780,
    48'h000004214c698,
    48'h00000423551b8,
    48'h000004214c490,
    48'h0000042355190,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c494,
    48'h000004214c69c,
    48'h0000040139544,
    48'h000004214c344,
    48'h000004013885c,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136514,
    48'h000004214c781,
    48'h000004214c599,
    48'h00000423551c8,
    48'h0000040136800,
    48'h0000040138f44,
    48'h00000423551c8,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h0000040022cc4,
    48'h0000040022de8,
    48'h0000040022ccc,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000004214c69c,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8018,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034baa,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000007b034ff4,
    48'h000004214c344,
    48'h000004013885c,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c344,
    48'h0000040139544,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h0000040021af0,
    48'h0000040021af8,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h0000040138eb0,
    48'h0000040138eb1,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h0000040138eb0,
    48'h0000040138eb1,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c780,
    48'h0000040139978,
    48'h000004214c490,
    48'h0000042355190,
    48'h0000040138f40,
    48'h0000042355190,
    48'h000004214c490,
    48'h0000040139978,
    48'h000004214c698,
    48'h0000042355190,
    48'h0000042355190,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c490,
    48'h0000040139540,
    48'h000007b035194,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355194,
    48'h0000042355190,
    48'h0000042355180,
    48'h00000400015bc,
    48'h00000423551e8,
    48'h0000042355150,
    48'h0000042355150,
    48'h000007b035154,
    48'h0000042355154,
    48'h000004213a120,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h0000042355148,
    48'h0000042355190,
    48'h0000042355130,
    48'h0000042355192,
    48'h0000042355132,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h0000042355194,
    48'h0000042355134,
    48'h0000042355180,
    48'h0000042355120,
    48'h0000042355182,
    48'h0000042355122,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h0000042355188,
    48'h0000042355128,
    48'h0000042355178,
    48'h0000042355118,
    48'h000004235517c,
    48'h000004235511c,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355158,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e8,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h00000423550c0,
    48'h0000042355048,
    48'h0000042355048,
    48'h000007b035154,
    48'h000004235504c,
    48'h000004213a120,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042355040,
    48'h0000042354d90,
    48'h000004235503c,
    48'h0000042355190,
    48'h0000042351df0,
    48'h0000042355050,
    48'h0000042355798,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040023890,
    48'h0000040023b38,
    48'h000007b034f11,
    48'h0000040139540,
    48'h0000040023b38,
    48'h00000400024b8,
    48'h0000040023b38,
    48'h0000040001fac,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040001fac,
    48'h0000040023b38,
    48'h000007b034f11,
    48'h0000040023b38,
    48'h0000040023a5a,
    48'h00000400237b0,
    48'h0000040023898,
    48'h0000040023b38,
    48'h000007b035158,
    48'h000007b03515c,
    48'h000007b035160,
    48'h000007b035164,
    48'h000007b035164,
    48'h000007b035160,
    48'h000004214c960,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b09e0,
    48'h00000423b09e0,
    48'h00000423b09e2,
    48'h0000040002104,
    48'h000004214c960,
    48'h0000000384108,
    48'h000007b03515c,
    48'h00000423b09e4,
    48'h000004214c960,
    48'h0000040023898,
    48'h0000040139978,
    48'h000007b034ff0,
    48'h0000040139978,
    48'h00000423b09e4,
    48'h00000401364c8,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000004214c344,
    48'h000004214c69c,
    48'h000004214c494,
    48'h000004013885c,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c781,
    48'h000004013997c,
    48'h000004214c494,
    48'h00000423551b8,
    48'h0000040138f44,
    48'h00000423551b8,
    48'h000004214c494,
    48'h000004013997c,
    48'h000004214c69c,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c494,
    48'h0000040139544,
    48'h000007b035194,
    48'h00000423551b8,
    48'h00000423551b8,
    48'h00000423551bc,
    48'h00000423551b8,
    48'h00000423551a8,
    48'h00000400015bc,
    48'h00000423551e8,
    48'h0000042355150,
    48'h0000042355150,
    48'h000007b035154,
    48'h0000042355154,
    48'h000004213a120,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h0000042355148,
    48'h00000423551b8,
    48'h0000042355130,
    48'h00000423551ba,
    48'h0000042355132,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h00000423551bc,
    48'h0000042355134,
    48'h00000423551a8,
    48'h0000042355120,
    48'h00000423551aa,
    48'h0000042355122,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h00000423551b0,
    48'h0000042355128,
    48'h00000423551a0,
    48'h0000042355118,
    48'h00000423551a4,
    48'h000004235511c,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355158,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e8,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h00000423550c0,
    48'h0000042355048,
    48'h0000042355048,
    48'h000007b035154,
    48'h000004235504c,
    48'h000004213a120,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042355040,
    48'h0000042354d90,
    48'h000004235503c,
    48'h00000423551b8,
    48'h0000042351df0,
    48'h0000042355050,
    48'h0000042355798,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h0000040139978,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000042355190,
    48'h0000040138f40,
    48'h0000042355190,
    48'h00000400237b0,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000007b034ff4,
    48'h000004214c69c,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000007b034fb8,
    48'h0000040139978,
    48'h0000042355192,
    48'h000004214c780,
    48'h0000042355190,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035194,
    48'h0000042355190,
    48'h0000042355190,
    48'h0000042355194,
    48'h0000042355190,
    48'h0000042355180,
    48'h00000400015bc,
    48'h00000423551e8,
    48'h0000042355150,
    48'h0000042355150,
    48'h000007b035154,
    48'h0000042355160,
    48'h0000042355140,
    48'h0000042355144,
    48'h0000042355138,
    48'h0000042355148,
    48'h0000042355190,
    48'h0000042355130,
    48'h0000042355192,
    48'h0000042355132,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h0000042355194,
    48'h0000042355134,
    48'h0000042355180,
    48'h0000042355120,
    48'h0000042355182,
    48'h0000042355122,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h0000042355188,
    48'h0000042355128,
    48'h0000042355178,
    48'h0000042355118,
    48'h000004235517c,
    48'h000004235511c,
    48'h0000042355148,
    48'h0000042355130,
    48'h0000042355158,
    48'h00000423550e0,
    48'h00000423550e0,
    48'h00000423550e8,
    48'h00000423550b8,
    48'h00000423550b8,
    48'h00000423550c0,
    48'h0000042355048,
    48'h0000042355048,
    48'h000007b035154,
    48'h0000042355058,
    48'h0000042355038,
    48'h000004235503c,
    48'h0000042351df0,
    48'h0000042355040,
    48'h0000042354d90,
    48'h000004235503c,
    48'h0000042355190,
    48'h0000042351df0,
    48'h0000042355050,
    48'h0000042355798,
    48'h00000423b09e2,
    48'h0000042355190,
    48'h0000042355192,
    48'h0000042355190,
    48'h00000400015a4,
    48'h0000042355190,
    48'h00000423b09e2,
    48'h000004213a240,
    48'h000004235914c,
    48'h0000000df7828,
    48'h000007b035258,
    48'h000007b03525c,
    48'h000007b035260,
    48'h000007b035264,
    48'h000007b035264,
    48'h000007b035260,
    48'h000004214c93c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b09e8,
    48'h00000423b09e8,
    48'h00000423b09ea,
    48'h00000400020e0,
    48'h000004214c93c,
    48'h00000003840fc,
    48'h000007b03525c,
    48'h00000423b09ec,
    48'h000004214c93c,
    48'h00000003840fd,
    48'h000007b035258,
    48'h00000423b09f0,
    48'h000004214c93c,
    48'h00000423b09e8,
    48'h000004214c90c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b09f8,
    48'h00000423b09f8,
    48'h00000423b0a0c,
    48'h00000423b0a10,
    48'h00000423b0a08,
    48'h00000423b0a14,
    48'h0000040002394,
    48'h0000040002394,
    48'h00000423b09fc,
    48'h00000423551e8,
    48'h00000423b0a04,
    48'h00000423b0a00,
    48'h00000423b0a00,
    48'h000004235515c,
    48'h00000423551e8,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040023978,
    48'h0000040136800,
    48'h000004214c494,
    48'h000007b034fb9,
    48'h000004013997c,
    48'h00000400015a4,
    48'h000007b034fb9,
    48'h000004214c69c,
    48'h000007b034ff4,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h00000423b09e2,
    48'h0000040022cc0,
    48'h0000040022cb8,
    48'h00000423551c4,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h000004013997c,
    48'h0000040022cc8,
    48'h0000040138eb1,
    48'h0000040022de8,
    48'h00000423551f0,
    48'h00000423551d0,
    48'h00000423551d4,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h00000423551fc,
    48'h00000423b03f2,
    48'h00000423b03f8,
    48'h00000423551e0,
    48'h00000423551e0,
    48'h000004213c310,
    48'h000004235525c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af264,
    48'h0000042355250,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355252,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355260,
    48'h0000042355240,
    48'h0000042355244,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235526c,
    48'h0000042355250,
    48'h0000042355250,
    48'h000004213c310,
    48'h0000042355294,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af264,
    48'h0000042355288,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235528a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355298,
    48'h0000042355278,
    48'h000004235527c,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h0000042354c72,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h0000040023760,
    48'h000007b034ca8,
    48'h00000423552a4,
    48'h0000042355288,
    48'h0000042355288,
    48'h000004213c310,
    48'h00000423552bc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af268,
    48'h00000423552b0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423552b2,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423552c0,
    48'h00000423552a8,
    48'h00000423552a8,
    48'h00000423552cc,
    48'h00000423b0412,
    48'h00000423b0418,
    48'h00000423552b0,
    48'h00000423552b0,
    48'h000004213c310,
    48'h00000423552fc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af268,
    48'h00000423552f0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423552f2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355300,
    48'h00000423552e0,
    48'h00000423552e4,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235530c,
    48'h00000423552f0,
    48'h00000423552f0,
    48'h000004213c310,
    48'h0000042355324,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af268,
    48'h0000042355318,
    48'h0000042355318,
    48'h0000042355318,
    48'h0000042355318,
    48'h000004213c310,
    48'h0000042355104,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af268,
    48'h00000423550f8,
    48'h00000423550f8,
    48'h00000423550f8,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h00000423550f8,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423553a4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af26c,
    48'h0000042355398,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235539a,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423553a8,
    48'h0000042355388,
    48'h000004235538c,
    48'h0000042355380,
    48'h0000042355384,
    48'h0000042355390,
    48'h0000042355378,
    48'h0000042355388,
    48'h0000042355388,
    48'h0000042355390,
    48'h0000042355378,
    48'h0000042355388,
    48'h000004214c8a8,
    48'h00000423553ac,
    48'h00000423553ac,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h00000423553ac,
    48'h00000423553a8,
    48'h00000423553ac,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h000004235538c,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042355390,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042355380,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042355384,
    48'h00000401367d0,
    48'h000007b0345c8,
    48'h0000040136428,
    48'h000007b034a48,
    48'h000004013893c,
    48'h0000042355378,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h000004235537a,
    48'h000004235537c,
    48'h0000042355368,
    48'h0000042355368,
    48'h0000042355368,
    48'h0000042355368,
    48'h0000042355368,
    48'h000004235536c,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042355370,
    48'h0000042355360,
    48'h0000042355364,
    48'h0000042355368,
    48'h0000042355370,
    48'h0000042355360,
    48'h000004235536c,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h0000042355390,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042355380,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042355380,
    48'h0000042355384,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042355380,
    48'h0000040138938,
    48'h0000042355382,
    48'h000007b034f58,
    48'h0000042355384,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042355378,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042355378,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042355378,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042355378,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000000df84e8,
    48'h0000042355378,
    48'h0000000df84e9,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h000004235538c,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042355390,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042355380,
    48'h0000042355380,
    48'h0000042355384,
    48'h0000042355380,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000042355378,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042355378,
    48'h0000042355378,
    48'h0000042355378,
    48'h000004235537a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042355390,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042355390,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034bac,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h00000423553a8,
    48'h0000042355388,
    48'h000004235538c,
    48'h0000042355380,
    48'h0000042355380,
    48'h0000042355380,
    48'h0000042355384,
    48'h0000042355382,
    48'h0000040001fac,
    48'h0000040023a68,
    48'h0000040023768,
    48'h000007b034e30,
    48'h0000040023760,
    48'h000007b034cc8,
    48'h00000423553b4,
    48'h0000042355398,
    48'h0000042355398,
    48'h000004213c310,
    48'h00000423553fc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af26c,
    48'h00000423553f0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423553f2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355400,
    48'h00000423553e0,
    48'h00000423553e4,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h000004235540c,
    48'h00000423b0422,
    48'h00000423b0428,
    48'h00000423553f0,
    48'h00000423553f0,
    48'h000004213c310,
    48'h000004235546c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af26c,
    48'h0000042355460,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355462,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355470,
    48'h0000042355450,
    48'h0000042355454,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235547c,
    48'h0000042355460,
    48'h0000042355460,
    48'h000004213c310,
    48'h00000423554e4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af26c,
    48'h00000423554d8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423554da,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423554e8,
    48'h00000423554c8,
    48'h00000423554cc,
    48'h0000042351df0,
    48'h00000423554c8,
    48'h00000423554c8,
    48'h00000423554d0,
    48'h00000423554b8,
    48'h00000423554c8,
    48'h000004214c8a8,
    48'h00000423554ec,
    48'h00000423554ec,
    48'h000007b03508c,
    48'h0000000dfcf58,
    48'h000007b035094,
    48'h0000000df7bf8,
    48'h000007b035094,
    48'h00000423554ec,
    48'h00000423554e8,
    48'h00000423554ec,
    48'h00000400025e4,
    48'h00000423554d0,
    48'h0000040139dd0,
    48'h00000423554bc,
    48'h0000040138938,
    48'h00000423554d0,
    48'h0000040139dd4,
    48'h00000423554c0,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df88e0,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9d80,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df88e4,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9d84,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df8444,
    48'h0000000df8445,
    48'h0000000df8446,
    48'h0000000df8447,
    48'h0000000df8448,
    48'h0000000df8449,
    48'h0000000df844a,
    48'h0000000df844b,
    48'h0000000df844c,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df8450,
    48'h0000000df8451,
    48'h0000000df8452,
    48'h0000000df8453,
    48'h0000000df8454,
    48'h0000000df8455,
    48'h0000000df8456,
    48'h0000000df8457,
    48'h0000000df8458,
    48'h0000040138938,
    48'h00000423554a8,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df8444,
    48'h0000040138938,
    48'h0000040139dd0,
    48'h00000423554aa,
    48'h00000423554ac,
    48'h0000042355498,
    48'h0000042355498,
    48'h0000042355498,
    48'h0000042355498,
    48'h0000042355498,
    48'h000004235549c,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000423554a0,
    48'h0000042355490,
    48'h0000042355494,
    48'h0000042355498,
    48'h00000423554a0,
    48'h0000042355490,
    48'h000004235549c,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd0,
    48'h00000423554bc,
    48'h0000040138938,
    48'h000007b035050,
    48'h000004013893c,
    48'h00000423554b0,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df8450,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423554a8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df8444,
    48'h0000000df8444,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h00000423554a8,
    48'h0000000df8445,
    48'h00000423554a8,
    48'h0000000df8446,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h0000000df8447,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h00000423554a8,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423554b0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8450,
    48'h0000000df8450,
    48'h000007b0350bc,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h0000000df8451,
    48'h000007b034f5c,
    48'h0000040139a98,
    48'h000007b034f5c,
    48'h00000423554b0,
    48'h0000000df8452,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423554b0,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423554a8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df8448,
    48'h0000000df8448,
    48'h000007b0350bc,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h0000000df8449,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h00000423554a8,
    48'h0000000df844a,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423554b0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8453,
    48'h0000000df8453,
    48'h00000423554b0,
    48'h00000423554b4,
    48'h0000000df8454,
    48'h00000423554b0,
    48'h0000000df8455,
    48'h000007b034f5c,
    48'h0000040139a98,
    48'h000007b034f5c,
    48'h00000423554b0,
    48'h0000000df8456,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423554b0,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423554a8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df844b,
    48'h0000000df844b,
    48'h00000423554a8,
    48'h000007b034f40,
    48'h00000423554ac,
    48'h0000042355498,
    48'h0000000df844c,
    48'h000007b034f28,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h000007b0350a4,
    48'h00000423554a8,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423554b0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8457,
    48'h0000000df8457,
    48'h00000423554b0,
    48'h0000000df8458,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h000007b0350a4,
    48'h00000423554b0,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b034fd4,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423554bc,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423554c0,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000004013893c,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h000004013893c,
    48'h00000423554b4,
    48'h000007b034fa4,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h000007b034fa0,
    48'h000007b035018,
    48'h000007b035018,
    48'h0000040138938,
    48'h000007b035018,
    48'h000007b034fa0,
    48'h000007b035154,
    48'h000007b035018,
    48'h000007b035068,
    48'h000007b035150,
    48'h000007b035018,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb17b,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd0,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554aa,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423554bc,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423554bc,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fb8,
    48'h000007b035001,
    48'h000007b034fd4,
    48'h000007b034fec,
    48'h000007b035009,
    48'h000007b034fec,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb17c,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b4,
    48'h0000040136800,
    48'h0000040139540,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040139540,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c494,
    48'h000004214c69c,
    48'h0000040139544,
    48'h000004214c344,
    48'h000004013885c,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040136514,
    48'h000004214c781,
    48'h000004214c599,
    48'h00000423554c0,
    48'h0000040136800,
    48'h0000040138f44,
    48'h00000423554c0,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h0000040022cc4,
    48'h0000040022de8,
    48'h0000040022ccc,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000004214c69c,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8018,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034bad,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000007b034ff4,
    48'h000004214c344,
    48'h000004013885c,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c344,
    48'h0000040139544,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h0000040021af0,
    48'h0000040021af8,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h0000040138eb0,
    48'h0000040138eb1,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h000007b034f4a,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h000007b034f48,
    48'h000007b034f4b,
    48'h000007b034f49,
    48'h000007b034f4b,
    48'h000007b034f49,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040021ae0,
    48'h000007b034f48,
    48'h000007b034f4a,
    48'h0000040138eb1,
    48'h0000040138eb0,
    48'h0000040021ae8,
    48'h0000040021ae8,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c344,
    48'h000004214c69c,
    48'h000004214c494,
    48'h000004013885c,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c781,
    48'h000004013997c,
    48'h000004214c494,
    48'h00000423554b0,
    48'h0000040138f44,
    48'h00000423554b0,
    48'h000004214c494,
    48'h000004013997c,
    48'h000004214c69c,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c494,
    48'h0000040139544,
    48'h000007b035194,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554b0,
    48'h00000423554e0,
    48'h0000042355460,
    48'h0000042355460,
    48'h0000042355468,
    48'h00000423553f0,
    48'h00000423553f0,
    48'h000007b035154,
    48'h00000423553f4,
    48'h000004213a120,
    48'h0000042355400,
    48'h00000423553e0,
    48'h00000423553e8,
    48'h00000423553d0,
    48'h00000423554b0,
    48'h00000423553f8,
    48'h0000042355398,
    48'h0000042355398,
    48'h000007b035154,
    48'h000004235539c,
    48'h000004213a120,
    48'h00000423553a8,
    48'h0000042355388,
    48'h0000042355390,
    48'h0000042355378,
    48'h00000423554b0,
    48'h00000423553a0,
    48'h00000423550f8,
    48'h000004013997c,
    48'h0000040138eb1,
    48'h0000040139544,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040023890,
    48'h0000040023b38,
    48'h000007b034f11,
    48'h0000040139544,
    48'h0000040023b38,
    48'h0000040002490,
    48'h0000040023b38,
    48'h0000040001fac,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040001fac,
    48'h0000040023b38,
    48'h000007b034f11,
    48'h0000040023b38,
    48'h0000040023a5a,
    48'h00000400237b0,
    48'h0000040023898,
    48'h00000423b09e2,
    48'h000004013997c,
    48'h000007b034ff4,
    48'h000004013997c,
    48'h00000423b09e4,
    48'h00000401364c8,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c780,
    48'h0000040139978,
    48'h000004214c490,
    48'h00000423554a8,
    48'h0000040138f40,
    48'h00000423554a8,
    48'h000004214c490,
    48'h0000040139978,
    48'h000004214c698,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h000007b035154,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000004214c490,
    48'h0000040139540,
    48'h000007b035194,
    48'h00000423554a8,
    48'h00000423554a8,
    48'h00000423554ac,
    48'h00000423554a8,
    48'h0000042355498,
    48'h00000400015bc,
    48'h00000423554e0,
    48'h0000042355460,
    48'h0000042355460,
    48'h0000042355468,
    48'h00000423553f0,
    48'h00000423553f0,
    48'h000007b035154,
    48'h00000423553f4,
    48'h000004213a120,
    48'h0000042355400,
    48'h00000423553e0,
    48'h00000423553e4,
    48'h0000042351df0,
    48'h00000423553e8,
    48'h00000423553d0,
    48'h00000423553f8,
    48'h0000042355398,
    48'h0000042355398,
    48'h000007b035154,
    48'h000004235539c,
    48'h000004213a120,
    48'h00000423553a8,
    48'h0000042355388,
    48'h000004235538c,
    48'h0000042355380,
    48'h0000042355390,
    48'h00000423554a8,
    48'h0000042355378,
    48'h00000423554aa,
    48'h000004235537a,
    48'h000004214c96c,
    48'h0000040002110,
    48'h0000000384130,
    48'h00000423554ac,
    48'h000004235537c,
    48'h0000042355498,
    48'h0000042355368,
    48'h000004235549a,
    48'h000004235536a,
    48'h000004214c988,
    48'h000004000212c,
    48'h00000003840fd,
    48'h00000423554a0,
    48'h0000042355370,
    48'h0000042355490,
    48'h0000042355360,
    48'h0000042355494,
    48'h0000042355364,
    48'h0000042355390,
    48'h0000042355378,
    48'h00000423553a0,
    48'h00000423550f8,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff4,
    48'h000004013997c,
    48'h000004214c69c,
    48'h000004214c494,
    48'h00000423554b0,
    48'h0000040138f44,
    48'h00000423554b0,
    48'h00000400237b0,
    48'h0000040136800,
    48'h000007b034f4a,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000007b034fb8,
    48'h0000040139978,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h000004214c494,
    48'h000007b034fb9,
    48'h000004013997c,
    48'h00000423554b2,
    48'h000004214c344,
    48'h000004214c781,
    48'h00000423554b0,
    48'h00000423b09e2,
    48'h00000423554b0,
    48'h00000423554b2,
    48'h00000423554b0,
    48'h00000400015a4,
    48'h00000423554b0,
    48'h00000423b09e2,
    48'h000004213a240,
    48'h000004235914c,
    48'h0000000df7828,
    48'h000007b035258,
    48'h000007b03525c,
    48'h000007b035260,
    48'h000007b035264,
    48'h000007b035264,
    48'h000007b035260,
    48'h000004214c93c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b0a18,
    48'h00000423b0a18,
    48'h00000423b0a1a,
    48'h00000400020e0,
    48'h000004214c93c,
    48'h00000003840fc,
    48'h000007b03525c,
    48'h00000423b0a1c,
    48'h000004214c93c,
    48'h00000003840fd,
    48'h000007b035258,
    48'h00000423b0a20,
    48'h000004214c93c,
    48'h00000423b0a18,
    48'h000004214c90c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b0a28,
    48'h00000423b0a28,
    48'h00000423b0a3c,
    48'h00000423b0a40,
    48'h00000423b0a38,
    48'h00000423b0a44,
    48'h0000040002394,
    48'h0000040002394,
    48'h00000423b0a2c,
    48'h00000423554e0,
    48'h00000423b0a34,
    48'h00000423b0a30,
    48'h00000423b0a30,
    48'h000004235546c,
    48'h00000423554e0,
    48'h00000400015a4,
    48'h000007b034fb9,
    48'h000004214c69c,
    48'h000007b034ff4,
    48'h0000040023978,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h000004013997c,
    48'h00000423b09e2,
    48'h0000040022ccc,
    48'h0000040022cc4,
    48'h00000423554c0,
    48'h0000040022de8,
    48'h00000423554e8,
    48'h00000423554c8,
    48'h00000423554cc,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h00000423554f4,
    48'h00000423554d8,
    48'h00000423554d8,
    48'h000004213c310,
    48'h0000042355554,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af270,
    48'h0000042355548,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235554a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355558,
    48'h0000042355538,
    48'h000004235553c,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042355564,
    48'h0000042355548,
    48'h0000042355548,
    48'h000004213c310,
    48'h000004235534c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af270,
    48'h0000042355340,
    48'h0000042355340,
    48'h0000042355340,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042355340,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423555e4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h00000423555d8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423555da,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423555e8,
    48'h00000423555c8,
    48'h00000423555cc,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h0000042354c72,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h0000040023760,
    48'h000007b034ca8,
    48'h00000423555f4,
    48'h00000423555d8,
    48'h00000423555d8,
    48'h000004213c310,
    48'h000004235560c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042355600,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355602,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355610,
    48'h00000423555f8,
    48'h00000423555f8,
    48'h000004235561c,
    48'h00000423b0442,
    48'h00000423b0448,
    48'h0000042355600,
    48'h0000042355600,
    48'h000004213c310,
    48'h000004235564c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042355640,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355642,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355650,
    48'h0000042355630,
    48'h0000042355634,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235565c,
    48'h0000042355640,
    48'h0000042355640,
    48'h000004213c310,
    48'h0000042355674,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042355668,
    48'h0000042355668,
    48'h0000042355668,
    48'h0000042355668,
    48'h000004213c310,
    48'h0000042355684,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042355678,
    48'h0000042355678,
    48'h0000042355678,
    48'h0000042355678,
    48'h000004213c310,
    48'h0000042354f84,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af274,
    48'h0000042354f78,
    48'h0000042354f78,
    48'h0000042354f78,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042354f78,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423556d4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h00000423556c8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423556ca,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423556d8,
    48'h00000423556b8,
    48'h00000423556bc,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000423556c0,
    48'h00000423556b0,
    48'h00000423556b8,
    48'h00000423556b8,
    48'h00000423556c0,
    48'h00000423556b0,
    48'h00000423556b8,
    48'h000004214c8a8,
    48'h00000423556dc,
    48'h00000423556dc,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h00000423556dc,
    48'h00000423556d8,
    48'h00000423556dc,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h00000423556bc,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h00000423556c0,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354d00,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040136428,
    48'h000007b034a54,
    48'h000004013893c,
    48'h00000423556b0,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h00000423556b2,
    48'h00000423556b4,
    48'h00000423556a0,
    48'h00000423556a0,
    48'h00000423556a0,
    48'h00000423556a0,
    48'h00000423556a0,
    48'h00000423556a4,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000423556a8,
    48'h0000042355698,
    48'h000004235569c,
    48'h00000423556a0,
    48'h00000423556a8,
    48'h0000042355698,
    48'h00000423556a4,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h00000401367d0,
    48'h000007b0345d4,
    48'h0000040139dd4,
    48'h00000423556c0,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042354d00,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042354d00,
    48'h0000040138938,
    48'h0000042354d02,
    48'h000007b034f58,
    48'h0000042354d04,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423556b0,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h00000423556b0,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h00000423556b0,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h00000423556b0,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h0000000df84e8,
    48'h00000423556b0,
    48'h0000000df84e9,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423556bc,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423556c0,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042354d00,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b0,
    48'h00000423556b2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423556c0,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423556c0,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034baf,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h00000423556d8,
    48'h00000423556b8,
    48'h00000423556bc,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d00,
    48'h0000042354d04,
    48'h0000042354d02,
    48'h0000040001fac,
    48'h0000040023a6e,
    48'h0000040023768,
    48'h000007b034e33,
    48'h0000040023760,
    48'h000007b034cd4,
    48'h00000423556e4,
    48'h00000423556c8,
    48'h00000423556c8,
    48'h000004213c310,
    48'h000004235572c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042355720,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355722,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h0000042355730,
    48'h0000042355710,
    48'h0000042355714,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042355718,
    48'h0000042355708,
    48'h0000042355710,
    48'h0000042355710,
    48'h0000042355718,
    48'h0000042355708,
    48'h0000042355710,
    48'h000004214c8a8,
    48'h0000042355734,
    48'h0000042355734,
    48'h000007b03508c,
    48'h0000000dfcfa8,
    48'h000007b035094,
    48'h0000000df7c48,
    48'h000007b035094,
    48'h0000042355734,
    48'h0000042355730,
    48'h0000042355734,
    48'h0000040002634,
    48'h0000040139dd0,
    48'h0000042355714,
    48'h0000040139dd4,
    48'h0000040138938,
    48'h0000042355718,
    48'h000004013893c,
    48'h000007b03508c,
    48'h0000000df8a70,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000df9f10,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df8a74,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000df9f14,
    48'h000007b03506c,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000000df84d5,
    48'h0000000df84d6,
    48'h0000000df84d7,
    48'h0000000df84d8,
    48'h0000000df84d9,
    48'h0000000df84da,
    48'h0000000df84db,
    48'h0000000df84dc,
    48'h0000000df84dd,
    48'h0000000df84de,
    48'h0000000df84df,
    48'h0000000df84e0,
    48'h0000000df84e1,
    48'h0000000df84e2,
    48'h0000000df84e3,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h0000000df84e5,
    48'h0000000df84e6,
    48'h0000000df84e7,
    48'h0000000df84e8,
    48'h0000000df84e9,
    48'h0000000df84ea,
    48'h0000000df84eb,
    48'h0000000df84ec,
    48'h0000000df84ed,
    48'h0000000df84ee,
    48'h0000000df84ef,
    48'h0000000df84f0,
    48'h0000000df84f1,
    48'h0000000df84f2,
    48'h0000000df84f3,
    48'h0000000df84f4,
    48'h0000000df84f5,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df84d4,
    48'h0000040138938,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040136428,
    48'h000007b034a50,
    48'h000004013893c,
    48'h0000042355708,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df84e4,
    48'h000004013893c,
    48'h0000040139dd4,
    48'h000004235570a,
    48'h000004235570c,
    48'h00000423556f8,
    48'h00000423556f8,
    48'h00000423556f8,
    48'h00000423556f8,
    48'h00000423556f8,
    48'h00000423556fc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042355700,
    48'h00000423556f0,
    48'h00000423556f4,
    48'h00000423556f8,
    48'h0000042355700,
    48'h00000423556f0,
    48'h00000423556fc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h00000401367d0,
    48'h000007b0345d0,
    48'h0000040139dd4,
    48'h0000042355718,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h0000042354d90,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df84d4,
    48'h0000000df84d4,
    48'h000007b035018,
    48'h0000000df84d5,
    48'h000007b0350bc,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h000007b034f58,
    48'h0000040139a98,
    48'h000007b034f58,
    48'h0000042354d90,
    48'h0000040138938,
    48'h0000042354d92,
    48'h000007b034f58,
    48'h0000042354d94,
    48'h00000400024b8,
    48'h0000040001fac,
    48'h0000000df84d6,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042355708,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df84e4,
    48'h0000000df84e4,
    48'h000007b034f5c,
    48'h0000040139a84,
    48'h000007b034f5c,
    48'h0000042355708,
    48'h0000000df84e5,
    48'h000007b034f5c,
    48'h0000040139bac,
    48'h000007b034f5c,
    48'h0000042355708,
    48'h0000000df84e6,
    48'h000007b034f5c,
    48'h00000401364c8,
    48'h0000040139ca0,
    48'h000007b034f5c,
    48'h0000042355708,
    48'h0000000df84e7,
    48'h000007b0350bc,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000000df84e8,
    48'h0000042355708,
    48'h0000000df84e9,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000000df84ea,
    48'h000007b034f2c,
    48'h000007b034f5c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b035000,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b035001,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b03509c,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b035000,
    48'h000007b035001,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h0000042355714,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h0000042355718,
    48'h000007b034fbc,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035000,
    48'h000007b034fe8,
    48'h000007b034fd0,
    48'h00000400015a4,
    48'h0000040138938,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d90,
    48'h000007b035001,
    48'h000007b034fec,
    48'h000007b034fd4,
    48'h00000400015a4,
    48'h000004013893c,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000042355708,
    48'h000007b034fa4,
    48'h000007b03501c,
    48'h000007b03501c,
    48'h000004013893c,
    48'h000007b03501c,
    48'h000007b034fa4,
    48'h000007b035154,
    48'h000007b03501c,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b03501c,
    48'h000007b03514c,
    48'h000007b03508c,
    48'h0000000dfb1e0,
    48'h000007b035148,
    48'h000007b035144,
    48'h0000040139dd4,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042355708,
    48'h0000042355708,
    48'h0000042355708,
    48'h000004235570a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h0000042355718,
    48'h0000040136800,
    48'h0000040138f40,
    48'h0000042355718,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h000007b034fbc,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h000007b03508c,
    48'h0000000df8068,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034baf,
    48'h0000040138eb0,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001f9c,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h000004214c490,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h0000040022cbc,
    48'h0000040138eb0,
    48'h0000040022de8,
    48'h0000042355730,
    48'h0000042355710,
    48'h0000042355714,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d90,
    48'h0000042354d94,
    48'h0000042354d92,
    48'h0000040001fac,
    48'h0000040023a6c,
    48'h0000040023768,
    48'h000007b034e32,
    48'h0000040023760,
    48'h000007b034cd0,
    48'h000004235573c,
    48'h0000042355720,
    48'h0000042355720,
    48'h000004213c310,
    48'h0000042355784,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042355778,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235577a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355788,
    48'h0000042355750,
    48'h0000042355754,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h0000040023a5e,
    48'h0000040023768,
    48'h000007b034e2b,
    48'h0000040023760,
    48'h000007b034cb4,
    48'h0000042355794,
    48'h0000042355778,
    48'h0000042355778,
    48'h000004213c310,
    48'h0000042354fac,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042354fa0,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042354fa2,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042354fb0,
    48'h0000042354f90,
    48'h0000042354f94,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042354fbc,
    48'h0000042354fa0,
    48'h0000042354fa0,
    48'h000004213c310,
    48'h000004235501c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042355010,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355012,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355020,
    48'h0000042355000,
    48'h0000042355004,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h000004235502c,
    48'h0000042355010,
    48'h0000042355010,
    48'h000004213c310,
    48'h000004235586c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h0000042355860,
    48'h0000042355860,
    48'h0000042355860,
    48'h0000042355860,
    48'h000004213c310,
    48'h00000423b034c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af278,
    48'h00000423b0340,
    48'h00000423b0340,
    48'h00000423b0340,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h00000423b0340,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h0000042354f54,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af27c,
    48'h0000042354f48,
    48'h0000042354f48,
    48'h0000042354f48,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042354f48,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423558c4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af280,
    48'h00000423558b8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423558ba,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423558c8,
    48'h00000423558a8,
    48'h00000423558ac,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h00000423558d4,
    48'h00000423b0462,
    48'h00000423b0468,
    48'h00000423558b8,
    48'h00000423558b8,
    48'h000004213c310,
    48'h0000042355934,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af280,
    48'h0000042355928,
    48'h0000040023768,
    48'h000004214c578,
    48'h000004235592a,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355938,
    48'h0000042355918,
    48'h000004235591c,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042355944,
    48'h0000042355928,
    48'h0000042355928,
    48'h000004213c310,
    48'h000004235596c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af280,
    48'h0000042355960,
    48'h0000040023768,
    48'h000004214c578,
    48'h0000042355962,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000042355970,
    48'h0000042355950,
    48'h0000042355954,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h0000042351df0,
    48'h000004235597c,
    48'h00000423b0472,
    48'h00000423b0478,
    48'h0000042355960,
    48'h0000042355960,
    48'h000004213c310,
    48'h00000423559dc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af284,
    48'h00000423559d0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423559d2,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423559e0,
    48'h00000423559c0,
    48'h00000423559c4,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h00000423559ec,
    48'h00000423559d0,
    48'h00000423559d0,
    48'h000004213c310,
    48'h000004235589c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af284,
    48'h0000042355890,
    48'h0000042355890,
    48'h0000042355890,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042355890,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423acd0c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h00000423acd00,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acd02,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423acd10,
    48'h00000423accf0,
    48'h00000423accf4,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c70,
    48'h0000042354c74,
    48'h0000042354c72,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h0000040023760,
    48'h000007b034ca8,
    48'h00000423acd1c,
    48'h00000423acd00,
    48'h00000423acd00,
    48'h000004213c310,
    48'h00000423acd34,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h00000423acd28,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acd2a,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423acd38,
    48'h00000423acd20,
    48'h00000423acd20,
    48'h00000423acd44,
    48'h00000423b0482,
    48'h00000423b0488,
    48'h00000423acd28,
    48'h00000423acd28,
    48'h000004213c310,
    48'h00000423acd74,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h00000423acd68,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acd6a,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423acd78,
    48'h00000423acd58,
    48'h00000423acd5c,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h0000042351de8,
    48'h00000423acd84,
    48'h00000423acd68,
    48'h00000423acd68,
    48'h000004213c310,
    48'h00000423acd9c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h00000423acd90,
    48'h00000423acd90,
    48'h00000423acd90,
    48'h00000423acd90,
    48'h000004213c310,
    48'h0000042355884,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af288,
    48'h0000042355878,
    48'h0000042355878,
    48'h0000042355878,
    48'h0000040023890,
    48'h00000400237b0,
    48'h0000040023890,
    48'h0000042355878,
    48'h0000040023890,
    48'h0000040023b38,
    48'h0000040136481,
    48'h00000400237b0,
    48'h0000040023890,
    48'h000004213c310,
    48'h00000423acde4,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423acdd8,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acdda,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423acde8,
    48'h00000423acdc8,
    48'h00000423acdcc,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h00000423acdd0,
    48'h00000423acdb8,
    48'h00000423acdc8,
    48'h00000423acdc8,
    48'h00000423acdd0,
    48'h00000423acdb8,
    48'h00000423acdc8,
    48'h000004214c8a8,
    48'h00000423acdec,
    48'h00000423acdec,
    48'h000007b03508c,
    48'h0000000dfd1c8,
    48'h000007b035094,
    48'h0000000df7e68,
    48'h000007b035094,
    48'h00000423acdec,
    48'h00000423acde8,
    48'h00000423acdec,
    48'h0000040002854,
    48'h0000040139dd0,
    48'h00000423acdcc,
    48'h0000040138938,
    48'h00000423acdd0,
    48'h0000040139dd4,
    48'h00000423acdbc,
    48'h000004013893c,
    48'h00000423acdd0,
    48'h0000040139dd8,
    48'h00000423acdc0,
    48'h0000040138940,
    48'h000007b03508c,
    48'h0000000df9510,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000dfa9b0,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df9514,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000dfa9b4,
    48'h000007b03506c,
    48'h000007b03508c,
    48'h0000000df9518,
    48'h000007b034f18,
    48'h000007b034f30,
    48'h0000000dfa9b8,
    48'h000007b035070,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df85f0,
    48'h0000000df85f1,
    48'h0000000df85f2,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df85f4,
    48'h0000040138938,
    48'h000004013893c,
    48'h00000423acdb0,
    48'h0000042354e20,
    48'h00000423acdb4,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h000007b035031,
    48'h0000000df85f5,
    48'h0000040138940,
    48'h000007b035058,
    48'h000007b034f30,
    48'h0000000df8750,
    48'h0000000df8751,
    48'h0000000df8752,
    48'h0000040138938,
    48'h00000423acdb0,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df85f0,
    48'h0000040138938,
    48'h00000423acdb4,
    48'h00000401367d0,
    48'h000007b0345a8,
    48'h0000040136428,
    48'h000007b034a28,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df85f4,
    48'h000004013893c,
    48'h0000042354e24,
    48'h00000401367d0,
    48'h000007b0345b4,
    48'h0000040136428,
    48'h000007b034a34,
    48'h0000040138940,
    48'h00000423acda8,
    48'h000007b035020,
    48'h000007b034f48,
    48'h000007b034f30,
    48'h0000000df8750,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acdb0,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df85f0,
    48'h0000000df85f0,
    48'h000007b035018,
    48'h0000000df85f1,
    48'h000007b034f58,
    48'h0000040139a84,
    48'h000007b034f58,
    48'h00000423acdb0,
    48'h0000040138938,
    48'h00000423acdb2,
    48'h000007b034f58,
    48'h00000423acdb4,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df85f2,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h0000042354e20,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df85f4,
    48'h0000000df85f4,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035031,
    48'h000007b034f70,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b034f58,
    48'h000007b035150,
    48'h000007b035154,
    48'h000004013893c,
    48'h0000040138938,
    48'h0000040139dd4,
    48'h0000040139dd0,
    48'h000007b035154,
    48'h000007b035150,
    48'h00000423acdb0,
    48'h0000042354e20,
    48'h00000423acdb2,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h0000040001fac,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h0000040139db0,
    48'h00000423acdbc,
    48'h0000040138950,
    48'h00000423afb50,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h0000040022e60,
    48'h00000423acde8,
    48'h00000423acdc8,
    48'h00000423acdcc,
    48'h00000423acdb0,
    48'h00000423acdd0,
    48'h00000423acdb8,
    48'h000004214c9c0,
    48'h0000040002164,
    48'h00000003840fd,
    48'h00000423acdc0,
    48'h00000423acda8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h00000003840fc,
    48'h00000423acdbc,
    48'h0000042351df8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h0000040002490,
    48'h00000423acdbc,
    48'h0000040022e70,
    48'h0000042354e20,
    48'h0000040022e60,
    48'h00000423acdb4,
    48'h00000423acdf4,
    48'h00000423b0522,
    48'h00000423b0524,
    48'h0000042354e24,
    48'h00000423b0528,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df85f5,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h0000042354e20,
    48'h000007b034f5c,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423acda8,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df8750,
    48'h0000000df8750,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423acda8,
    48'h0000000df8751,
    48'h00000423acda8,
    48'h00000423acdac,
    48'h0000000df8752,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b0350bc,
    48'h000007b034f72,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b034f60,
    48'h000007b034fa8,
    48'h000007b034f72,
    48'h000007b035002,
    48'h000007b034f7a,
    48'h000007b03500a,
    48'h000007b034f90,
    48'h000007b034fd8,
    48'h000007b034f82,
    48'h000007b035012,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b034ff0,
    48'h000007b035000,
    48'h000007b034fd0,
    48'h000007b035001,
    48'h000007b034fd4,
    48'h000007b034fe8,
    48'h000007b035002,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423acdcc,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423acdbc,
    48'h000007b034fbc,
    48'h0000040139dd8,
    48'h000007b035058,
    48'h00000423acdc0,
    48'h000007b034fc0,
    48'h000007b035000,
    48'h0000040138938,
    48'h00000423acdb0,
    48'h00000423acdb0,
    48'h000007b035001,
    48'h000004013893c,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h000007b035002,
    48'h000007b035000,
    48'h000007b034fd0,
    48'h000007b034fe8,
    48'h000007b035018,
    48'h000007b035018,
    48'h000007b034fe8,
    48'h000007b03501c,
    48'h000007b034fa0,
    48'h000007b035154,
    48'h000007b034fe8,
    48'h000007b03506c,
    48'h000007b035150,
    48'h000007b035068,
    48'h000007b035148,
    48'h000007b035144,
    48'h000007b03514c,
    48'h000004013893c,
    48'h0000040138938,
    48'h0000040139dd4,
    48'h0000040139dd0,
    48'h000007b035150,
    48'h000007b03514c,
    48'h000007b035148,
    48'h000007b035154,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h0000042354e20,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h0000042354e20,
    48'h0000042354e22,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000004214c698,
    48'h0000040139540,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040139978,
    48'h0000040138eb0,
    48'h0000040136510,
    48'h000004214c780,
    48'h000004214c598,
    48'h00000423acdbc,
    48'h0000040136800,
    48'h0000040138f40,
    48'h00000423acdbc,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040022cb8,
    48'h0000040022de8,
    48'h0000040022cc0,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h0000040022cc4,
    48'h0000040022de8,
    48'h0000040022ccc,
    48'h0000040139978,
    48'h0000040139540,
    48'h000007b035210,
    48'h000007b035214,
    48'h000007b035214,
    48'h000007b035210,
    48'h00000423acdb0,
    48'h0000042354e20,
    48'h00000423acdb2,
    48'h0000042354e22,
    48'h0000040001fac,
    48'h0000040001fac,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h0000040139db0,
    48'h00000423acdbc,
    48'h0000040138950,
    48'h00000423afb50,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h0000040022e60,
    48'h00000423acde8,
    48'h00000423acdc8,
    48'h00000423acdcc,
    48'h00000423acdb0,
    48'h00000423acdd0,
    48'h00000423acdb8,
    48'h000004214c9c0,
    48'h0000040002164,
    48'h00000003840fd,
    48'h00000423acdc0,
    48'h00000423acda8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h00000003840fc,
    48'h00000423acdbc,
    48'h0000042351df8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h0000040002490,
    48'h00000423acdbc,
    48'h0000040022e70,
    48'h0000042354e20,
    48'h0000040022e60,
    48'h00000423acdb4,
    48'h00000423acdf4,
    48'h00000423b0522,
    48'h00000423b0524,
    48'h0000042354e24,
    48'h00000423b0528,
    48'h0000040139978,
    48'h0000042354e20,
    48'h000007b03520c,
    48'h000007b035210,
    48'h0000040022e78,
    48'h000007b035214,
    48'h0000040022e60,
    48'h00000423acdb4,
    48'h000007b035254,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423acde0,
    48'h0000042355878,
    48'h0000040022e88,
    48'h000007b034fe8,
    48'h000007b034fbc,
    48'h0000040022e88,
    48'h000007b034fb8,
    48'h000007b035001,
    48'h000007b034fd4,
    48'h000007b035002,
    48'h000007b034ff0,
    48'h000007b034fd8,
    48'h00000400015a4,
    48'h0000040138940,
    48'h00000423acda8,
    48'h00000423acda8,
    48'h00000423acda8,
    48'h0000040136800,
    48'h000004214c698,
    48'h0000040136800,
    48'h0000040138eb0,
    48'h000004214c490,
    48'h000007b03508c,
    48'h0000000df8288,
    48'h0000040136800,
    48'h000004213c310,
    48'h000007b034bb4,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c340,
    48'h0000040138858,
    48'h0000040001fac,
    48'h0000040001fac,
    48'h000004214c340,
    48'h0000040139540,
    48'h0000040001fac,
    48'h0000040136800,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000004214c340,
    48'h000004214c698,
    48'h0000040138858,
    48'h0000040001fac,
    48'h0000040001fac,
    48'h000004214c780,
    48'h0000040139978,
    48'h0000040136800,
    48'h0000040136800,
    48'h000007b034f48,
    48'h000007b034ff0,
    48'h000004214c698,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h0000040023760,
    48'h0000040023768,
    48'h000007b034ca8,
    48'h000007b034e28,
    48'h0000040136800,
    48'h0000040136800,
    48'h000004214c490,
    48'h000007b034fb8,
    48'h0000040139978,
    48'h0000042354e22,
    48'h000004214c780,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423acdb2,
    48'h0000042354e20,
    48'h0000042354e22,
    48'h0000042354e20,
    48'h00000400015a4,
    48'h0000042354e20,
    48'h0000042354e24,
    48'h00000423acdb2,
    48'h000004213a240,
    48'h000004235914c,
    48'h0000000df7828,
    48'h000007b035258,
    48'h000007b03525c,
    48'h000007b035260,
    48'h000007b035264,
    48'h000007b035264,
    48'h000007b035260,
    48'h000004214c93c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b0a48,
    48'h00000423b0a48,
    48'h00000423b0a4a,
    48'h00000400020e0,
    48'h000004214c93c,
    48'h00000003840fc,
    48'h000007b03525c,
    48'h00000423b0a4c,
    48'h000004214c93c,
    48'h00000003840fd,
    48'h000007b035258,
    48'h00000423b0a50,
    48'h000004214c93c,
    48'h00000423b0a48,
    48'h000004214c90c,
    48'h000004213c320,
    48'h000004214c844,
    48'h000004214c848,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c844,
    48'h000004214c850,
    48'h000004214c844,
    48'h000004214c83c,
    48'h000004214c848,
    48'h000004214c840,
    48'h000004214c844,
    48'h000004214c840,
    48'h00000423b0a58,
    48'h00000423b0a58,
    48'h00000423b0a6c,
    48'h00000423b0a70,
    48'h00000423b0a68,
    48'h00000423b0a74,
    48'h0000040002394,
    48'h0000040002394,
    48'h00000423b0a5c,
    48'h00000423acde0,
    48'h00000423b0a64,
    48'h00000423b0a60,
    48'h00000423b0a60,
    48'h0000042355884,
    48'h00000423acde0,
    48'h00000400015a4,
    48'h000007b034fb8,
    48'h000004214c698,
    48'h0000040139978,
    48'h000007b034ff0,
    48'h0000040136800,
    48'h0000040022de8,
    48'h0000040022cbc,
    48'h0000040139978,
    48'h00000423acdb2,
    48'h0000040022cc0,
    48'h0000040022cb8,
    48'h00000423acdbc,
    48'h0000040022de8,
    48'h0000040022cc8,
    48'h0000040139978,
    48'h00000423acdb2,
    48'h0000040022ccc,
    48'h0000040022cc4,
    48'h00000423acdcc,
    48'h0000040022de8,
    48'h00000423acde8,
    48'h00000423acdc8,
    48'h00000423acdcc,
    48'h00000423acdb0,
    48'h00000423acdb0,
    48'h00000423acdb0,
    48'h00000423acdb4,
    48'h00000423acdb2,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h00000423acdf4,
    48'h00000423b0522,
    48'h00000423b0528,
    48'h00000423acdd8,
    48'h00000423acdd8,
    48'h000004213c310,
    48'h00000423ace24,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423ace18,
    48'h00000423ace18,
    48'h00000423ace18,
    48'h00000423ace18,
    48'h000004213c310,
    48'h00000423ace6c,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423ace60,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423ace62,
    48'h0000040136800,
    48'h0000040136800,
    48'h00000423ace70,
    48'h00000423ace50,
    48'h00000423ace54,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h00000423ace3c,
    48'h00000423ace3a,
    48'h0000040001fac,
    48'h0000040023a58,
    48'h0000040023768,
    48'h000007b034e28,
    48'h0000040023760,
    48'h000007b034ca8,
    48'h00000423ace7c,
    48'h00000423b0502,
    48'h00000423b0508,
    48'h00000423ace60,
    48'h00000423ace60,
    48'h000004213c310,
    48'h00000423aceac,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423acea0,
    48'h00000423acea0,
    48'h00000423acea0,
    48'h00000423acea0,
    48'h000004213c310,
    48'h00000423acefc,
    48'h0000040139620,
    48'h0000040139a58,
    48'h00000423af28c,
    48'h00000423acef0,
    48'h0000040023768,
    48'h000004214c578,
    48'h00000423acef2,
    48'h0000040023c88,
    48'h000007b034ed4,
    48'h000007b035084,
    48'h0000040036348,
    48'h0000040022e58,
    48'h0000040022cb0,
    48'h0000040022de8,
    48'h0000040022e68,
    48'h0000040136800,
    48'h0000040022e70,
    48'h0000040022e60,
    48'h000007b034ed4,
    48'h0000040022e78,
    48'h00000423acf00,
    48'h00000423acee0,
    48'h00000423acee4,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h00000423acee8,
    48'h00000423b0860,
    48'h00000423acee0,
    48'h00000423acee0,
    48'h00000423acee8,
    48'h00000423b0860,
    48'h00000423acee0,
    48'h000004214c8a8,
    48'h00000423acf04,
    48'h00000423acf04,
    48'h000007b03508c,
    48'h0000000dfd13c,
    48'h000007b035094,
    48'h0000000df7ddc,
    48'h000007b035094,
    48'h00000423acf04,
    48'h00000423acf00,
    48'h00000423acf04,
    48'h00000400027c8,
    48'h0000040139dd0,
    48'h00000423acee4,
    48'h0000040138938,
    48'h00000423acee8,
    48'h0000040139dd4,
    48'h00000423b0864,
    48'h000004013893c,
    48'h00000423acee8,
    48'h0000040139dd8,
    48'h00000423b0868,
    48'h0000040138940,
    48'h000007b03508c,
    48'h0000000df9254,
    48'h000007b034f10,
    48'h000007b034f28,
    48'h0000000dfa6f4,
    48'h000007b035068,
    48'h000007b03508c,
    48'h0000000df9258,
    48'h000007b034f14,
    48'h000007b034f2c,
    48'h0000000dfa6f8,
    48'h000007b03506c,
    48'h000007b03508c,
    48'h0000000df925c,
    48'h000007b034f18,
    48'h000007b034f30,
    48'h0000000dfa6fc,
    48'h000007b035070,
    48'h0000040138938,
    48'h000007b035050,
    48'h000007b034f28,
    48'h0000000df868c,
    48'h0000000df868d,
    48'h0000000df868e,
    48'h0000000df868f,
    48'h0000000df8690,
    48'h000004013893c,
    48'h000007b035054,
    48'h000007b034f2c,
    48'h0000000df8674,
    48'h0000000df8675,
    48'h0000040138938,
    48'h000004013893c,
    48'h00000423acec8,
    48'h00000423ace38,
    48'h00000423acecc,
    48'h00000423ace38,
    48'h00000423ace3c,
    48'h000007b035031,
    48'h0000040138938,
    48'h0000040138940,
    48'h00000423acec8,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h000007b035032,
    48'h0000000df8676,
    48'h0000000df8677,
    48'h0000040138938,
    48'h000004013893c,
    48'h00000423acec8,
    48'h00000423ace38,
    48'h00000423acecc,
    48'h00000423ace38,
    48'h00000423ace3c,
    48'h000007b035031,
    48'h0000040138938,
    48'h0000040138940,
    48'h00000423acec8,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h000007b035032,
    48'h0000000df8678,
    48'h0000040138940,
    48'h000007b035058,
    48'h000007b034f30,
    48'h0000000df8728,
    48'h0000000df8729,
    48'h0000000df872a,
    48'h0000000df872b,
    48'h0000000df872c,
    48'h0000000df872d,
    48'h0000000df872e,
    48'h0000000df872f,
    48'h0000000df8730,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b035018,
    48'h000007b034f40,
    48'h000007b034f28,
    48'h0000000df868c,
    48'h0000040138938,
    48'h00000423acecc,
    48'h00000401367d0,
    48'h000007b0345a8,
    48'h0000040136428,
    48'h000007b034a28,
    48'h000004013893c,
    48'h00000423ace38,
    48'h000007b03501c,
    48'h000007b034f44,
    48'h000007b034f2c,
    48'h0000000df8674,
    48'h000004013893c,
    48'h00000423ace3c,
    48'h00000401367d0,
    48'h000007b0345a8,
    48'h0000040136428,
    48'h000007b034a28,
    48'h0000040138940,
    48'h00000423b0848,
    48'h000007b035020,
    48'h000007b034f48,
    48'h000007b034f30,
    48'h0000000df8728,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df868c,
    48'h0000000df868c,
    48'h000007b035018,
    48'h0000000df868d,
    48'h000007b0350bc,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h00000423acec8,
    48'h00000423acec8,
    48'h0000000df868e,
    48'h000007b034f28,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h000007b0350a4,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f88,
    48'h000007b0350a4,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423ace38,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8674,
    48'h0000000df8674,
    48'h0000000df8675,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035031,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df8676,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423ace38,
    48'h000007b034f5c,
    48'h000007b034f8c,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423b0848,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df8728,
    48'h0000000df8728,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423b0848,
    48'h0000000df8729,
    48'h00000423b0848,
    48'h00000423b084c,
    48'h0000000df872a,
    48'h00000423b0848,
    48'h0000000df872b,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b034f7a,
    48'h00000423b0848,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df868f,
    48'h0000000df868f,
    48'h000007b034f58,
    48'h0000040139a84,
    48'h000007b034f58,
    48'h00000423acec8,
    48'h0000040138938,
    48'h00000423aceca,
    48'h000007b034f58,
    48'h00000423acecc,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df8690,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423ace38,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8677,
    48'h0000000df8677,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035031,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df8678,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b0350bc,
    48'h000007b034f71,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423b0848,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df872c,
    48'h0000000df872c,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423b0848,
    48'h0000000df872d,
    48'h000007b0350bc,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h00000423b0848,
    48'h0000000df872e,
    48'h00000423b0848,
    48'h00000423b084c,
    48'h0000000df872f,
    48'h00000423b0848,
    48'h0000000df8730,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b034f7a,
    48'h00000423b0848,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b034fa0,
    48'h000007b034f70,
    48'h000007b035000,
    48'h000007b034f78,
    48'h000007b035008,
    48'h000007b034f88,
    48'h000007b034fd0,
    48'h000007b034f80,
    48'h000007b035010,
    48'h000007b034f5c,
    48'h000007b034fa4,
    48'h000007b034f71,
    48'h000007b035001,
    48'h000007b034f79,
    48'h000007b035009,
    48'h000007b034f8c,
    48'h000007b034fd4,
    48'h000007b034f81,
    48'h000007b035011,
    48'h000007b034f60,
    48'h000007b034fa8,
    48'h000007b034f72,
    48'h000007b035002,
    48'h000007b034f7a,
    48'h000007b03500a,
    48'h000007b034f90,
    48'h000007b034fd8,
    48'h000007b034f82,
    48'h000007b035012,
    48'h000007b03509c,
    48'h000007b035094,
    48'h000007b03509c,
    48'h000007b03509c,
    48'h000007b035058,
    48'h000004013893c,
    48'h000007b035054,
    48'h0000040138940,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df868c,
    48'h0000000df868c,
    48'h000007b035018,
    48'h0000000df868d,
    48'h000007b0350bc,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h00000423acec8,
    48'h00000423acec8,
    48'h0000000df868e,
    48'h000007b034f28,
    48'h000007b034f80,
    48'h000007b034f78,
    48'h000007b0350a4,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f88,
    48'h000007b0350a4,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423b0848,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8674,
    48'h0000000df8674,
    48'h0000000df8675,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035032,
    48'h000007b034f70,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b0350a4,
    48'h000007b034f58,
    48'h000007b035150,
    48'h000007b035154,
    48'h000004013893c,
    48'h0000040138938,
    48'h0000040139dd4,
    48'h0000040139dd0,
    48'h000007b035154,
    48'h000007b035150,
    48'h00000423acec8,
    48'h00000423b0848,
    48'h00000423aceca,
    48'h00000423b084a,
    48'h0000040001fac,
    48'h0000040001f9c,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h0000040139db0,
    48'h00000423b0864,
    48'h0000040138950,
    48'h00000423afb50,
    48'h00000423aceca,
    48'h0000040001fac,
    48'h0000040022e60,
    48'h00000423acf00,
    48'h00000423acee0,
    48'h00000423acee4,
    48'h00000423acec8,
    48'h00000423acee8,
    48'h00000423b0860,
    48'h000004214c9ac,
    48'h0000040002150,
    48'h00000003840fd,
    48'h00000423b0868,
    48'h00000423b0848,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h00000003840fc,
    48'h00000423b0864,
    48'h0000042351df8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h0000040002468,
    48'h00000423b0864,
    48'h0000040022e70,
    48'h00000423b0848,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df8676,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423b0848,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423ace38,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df8728,
    48'h0000000df8728,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423ace38,
    48'h0000040138940,
    48'h00000423ace3a,
    48'h000007b034f60,
    48'h00000423ace3c,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df8729,
    48'h00000423ace38,
    48'h0000000df872a,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h0000000df872b,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b0350bc,
    48'h000007b034f72,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b0350a4,
    48'h000007b0350ac,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f28,
    48'h0000040138938,
    48'h00000423acec8,
    48'h000007b034f58,
    48'h000007b034f70,
    48'h000007b034f78,
    48'h000007b034f80,
    48'h000007b034f88,
    48'h0000000df868f,
    48'h0000000df868f,
    48'h000007b034f58,
    48'h0000040139a84,
    48'h000007b034f58,
    48'h00000423acec8,
    48'h0000040138938,
    48'h00000423aceca,
    48'h000007b034f58,
    48'h00000423acecc,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df8690,
    48'h000007b034f28,
    48'h000007b034f58,
    48'h000007b034f80,
    48'h000007b0350bc,
    48'h000007b034f70,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f2c,
    48'h000004013893c,
    48'h00000423b0848,
    48'h000007b034f5c,
    48'h000007b034f71,
    48'h000007b034f79,
    48'h000007b034f81,
    48'h000007b034f8c,
    48'h0000000df8677,
    48'h0000000df8677,
    48'h000007b034f8c,
    48'h000007b03509c,
    48'h000007b035032,
    48'h000007b034f70,
    48'h000007b034f70,
    48'h000007b034f58,
    48'h000007b034f58,
    48'h000007b035150,
    48'h000007b035154,
    48'h000004013893c,
    48'h0000040138938,
    48'h0000040139dd4,
    48'h0000040139dd0,
    48'h000007b035154,
    48'h000007b035150,
    48'h00000423acec8,
    48'h00000423b0848,
    48'h00000423aceca,
    48'h00000423b084a,
    48'h0000040001fac,
    48'h0000040001f9c,
    48'h00000423acec8,
    48'h00000423acecc,
    48'h0000040139db0,
    48'h00000423b0864,
    48'h0000040138950,
    48'h00000423afb50,
    48'h00000423aceca,
    48'h0000040001fac,
    48'h0000040022e60,
    48'h00000423acf00,
    48'h00000423acee0,
    48'h00000423acee4,
    48'h00000423acec8,
    48'h00000423acee8,
    48'h00000423b0860,
    48'h000004214c9ac,
    48'h0000040002150,
    48'h00000003840fd,
    48'h00000423b0868,
    48'h00000423b0848,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h00000003840fc,
    48'h00000423b0864,
    48'h0000042351df8,
    48'h000004214c950,
    48'h00000400020f4,
    48'h0000000384108,
    48'h0000000384108,
    48'h0000040002490,
    48'h00000423b0864,
    48'h0000040022e70,
    48'h00000423b0848,
    48'h000007b034f58,
    48'h000007b034f5c,
    48'h0000000df8678,
    48'h000007b034f2c,
    48'h000007b034f81,
    48'h000007b034f79,
    48'h00000423b0848,
    48'h000007b0350bc,
    48'h000007b0350b4,
    48'h000007b034f30,
    48'h0000040138940,
    48'h00000423ace38,
    48'h000007b034f60,
    48'h000007b034f72,
    48'h000007b034f7a,
    48'h000007b034f82,
    48'h000007b034f90,
    48'h0000000df872c,
    48'h0000000df872c,
    48'h000007b034f60,
    48'h0000040139a84,
    48'h000007b034f60,
    48'h00000423ace38,
    48'h0000040138940,
    48'h00000423ace3a,
    48'h000007b034f60,
    48'h00000423ace3c,
    48'h0000040002490,
    48'h0000040001fac,
    48'h0000000df872d,
    48'h000007b0350bc,
    48'h00000423ace38,
    48'h00000423ace3c,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h0000000df872e,
    48'h00000423ace38,
    48'h0000000df872f,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h00000423ace38,
    48'h0000000df8730,
    48'h000007b034f30,
    48'h000007b034f60,
    48'h000007b034f82,
    48'h000007b0350bc,
    48'h000007b034f72,
    48'h000007b034f80,
    48'h000007b034f81,
    48'h000007b034f82,
    48'h000007b0350ac,
    48'h000007b0350a4,
    48'h000007b035094,
    48'h000007b03509c,
    48'h000007b03509c,
    48'h000007b035054,
    48'h000004013893c,
    48'h000007b035058,
    48'h0000040138940,
    48'h000007b034fe8,
    48'h000007b034fec,
    48'h000007b034ff0,
    48'h000007b035000,
    48'h000007b035001,
    48'h000007b035002,
    48'h000007b034fd8,
    48'h0000040139dd0,
    48'h000007b035050,
    48'h00000423acee4,
    48'h000007b034fb8,
    48'h0000040139dd4,
    48'h000007b035054,
    48'h00000423b0864,
    48'h000007b034fbc,
    48'h0000040139dd8,
    48'h000007b035058
    };
endmodule
