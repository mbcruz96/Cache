
parameter SIZE = 1000;
module trace_addr(
    reg[31:0] test_addrs[0:SIZE-1]);
    
    assign test_addrs = 
    {
        48'h0000040020760,
        48'h000007b0337fc,
        48'h000007b0345f4,
        48'h000007b0337fc,
        48'h0000040059770,
        48'h000007b034514,
        48'h0000040059770,
        48'h0000040020464,
        48'h000007b0337fc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034514,
        48'h00000400ed7b4,
        48'h00000400ed7b8,
        48'h000007b034400,
        48'h0000040020468,
        48'h000007b03454c,
        48'h000007b034548,
        48'h000007b03454c,
        48'h000007b034548,
        48'h0000040020500,
        48'h00000400321ec,
        48'h000004003bfb0,
        48'h0000040020500,
        48'h00000400321ec,
        48'h000004003bfb0,
        48'h00000400ed7c0,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c18,
        48'h0000040045c18,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034538,
        48'h000007b0337fc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000004002060c,
        48'h0000040020344,
        48'h000007b03448c,
        48'h000007b03448c,
        48'h000007b0344fc,
        48'h0000040020608,
        48'h000004002060c,
        48'h000004000e43c,
        48'h000007b0344fc,
        48'h000007b0344fc,
        48'h0000040059918,
        48'h000007b0337fc,
        48'h000007b0344fc,
        48'h00000400597c0,
        48'h0000040020608,
        48'h000007b03450c,
        48'h000007b034508,
        48'h000007b034504,
        48'h000007b03450c,
        48'h000007b034508,
        48'h000007b034504,
        48'h000007b0345b0,
        48'h000007b0345ac,
        48'h000007b0345a8,
        48'h000004002060c,
        48'h000004000e43c,
        48'h000007b0345b4,
        48'h000007b0345b4,
        48'h0000040059914,
        48'h00000400d602c,
        48'h000007b0345b0,
        48'h000007b0337fc,
        48'h000007b0345b0,
        48'h00000400e5434,
        48'h00000400e5438,
        48'h000007b0345ac,
        48'h000007b0345cc,
        48'h000007b0345cc,
        48'h0000040020530,
        48'h0000040020504,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032344,
        48'h000007b0345a8,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h000007b0345b0,
        48'h00000400e53e4,
        48'h000007b0337fc,
        48'h000007b0345b0,
        48'h00000400e5408,
        48'h000007b0345cc,
        48'h000007b0345c8,
        48'h000007b0345cc,
        48'h000007b0345c8,
        48'h000007b03463c,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003232c,
        48'h00000400e70c0,
        48'h000007b03464c,
        48'h000007b034648,
        48'h000007b034644,
        48'h000007b03464c,
        48'h000007b034648,
        48'h000007b034644,
        48'h000007b0337fc,
        48'h000007b03463c,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045bfc,
        48'h00000400321e8,
        48'h000004003232c,
        48'h00000400e70bc,
        48'h00000400e70c4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003232c,
        48'h00000400e70d8,
        48'h00000400e70d8,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0345b0,
        48'h00000400e53e0,
        48'h000007b0345a8,
        48'h000007b034400,
        48'h00000400ed790,
        48'h000007b034404,
        48'h00000400ed794,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000004002078c,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034400,
        48'h000007b03440c,
        48'h000007b03440c,
        48'h0000040020530,
        48'h0000040020504,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032348,
        48'h0000040020628,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h00000400207bc,
        48'h000004002079c,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b03438c,
        48'h000007b03438c,
        48'h000007b03440c,
        48'h000007b03440c,
        48'h000007b03447c,
        48'h000004002078c,
        48'h0000040020610,
        48'h000007b0337fc,
        48'h0000040020614,
        48'h000004000e43c,
        48'h000007b03447c,
        48'h000007b03448c,
        48'h000007b03448c,
        48'h000007b03453c,
        48'h000007b034538,
        48'h000007b034534,
        48'h0000040020610,
        48'h0000040020614,
        48'h000004000e43c,
        48'h000007b03453c,
        48'h000007b03453c,
        48'h0000040059918,
        48'h000007b0337fc,
        48'h0000040020610,
        48'h00000400e5434,
        48'h00000400e53e8,
        48'h000007b03453c,
        48'h000007b03454c,
        48'h000007b034548,
        48'h000007b034544,
        48'h000007b034540,
        48'h000007b03454c,
        48'h000007b034548,
        48'h000007b034544,
        48'h000007b034540,
        48'h000007b0345fc,
        48'h000007b0345f8,
        48'h000007b0345f4,
        48'h000007b0345f0,
        48'h0000040020748,
        48'h000007b0345ec,
        48'h0000040058f58,
        48'h000007b0345ec,
        48'h000007b0345e8,
        48'h000007b034538,
        48'h00000400e5400,
        48'h000007b03460c,
        48'h000007b034608,
        48'h000007b03460c,
        48'h000007b034608,
        48'h000007b03468c,
        48'h000007b034688,
        48'h000007b03468c,
        48'h000007b034688,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045bf4,
        48'h00000400321e8,
        48'h0000040032324,
        48'h00000400e6aac,
        48'h00000400e6ab4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032324,
        48'h00000400e6acc,
        48'h000007b034534,
        48'h00000400e6acc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034534,
        48'h00000400e5404,
        48'h000007b03460c,
        48'h000007b034608,
        48'h000007b03460c,
        48'h000007b034608,
        48'h000007b03468c,
        48'h000007b034688,
        48'h000007b03468c,
        48'h000007b034688,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045bf8,
        48'h00000400321e8,
        48'h0000040032328,
        48'h00000400e6db4,
        48'h00000400e6dbc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032328,
        48'h00000400e6dd4,
        48'h000007b0345f8,
        48'h00000400e6dd4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0345f8,
        48'h000007b0337fc,
        48'h00000400e5418,
        48'h000007b03460c,
        48'h000007b034608,
        48'h000007b03460c,
        48'h000007b034608,
        48'h000007b03468c,
        48'h000007b034688,
        48'h000007b03468c,
        48'h000007b034688,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045bec,
        48'h00000400321e8,
        48'h000004003231c,
        48'h00000400e649c,
        48'h00000400e64a4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003231c,
        48'h00000400e64bc,
        48'h000007b0345fc,
        48'h00000400e64bc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0345fc,
        48'h000007b03460c,
        48'h000007b034608,
        48'h000007b034604,
        48'h000007b034600,
        48'h000007b03460c,
        48'h000007b034608,
        48'h000007b034604,
        48'h000007b034600,
        48'h000007b034694,
        48'h000007b034690,
        48'h000007b03468c,
        48'h000007b034688,
        48'h000007b034684,
        48'h0000040059770,
        48'h000007b034698,
        48'h0000040059774,
        48'h000007b03469c,
        48'h0000040059778,
        48'h000007b0346a0,
        48'h000004005977c,
        48'h000007b0346a4,
        48'h0000040059780,
        48'h000007b0346a8,
        48'h0000040059784,
        48'h000007b0346ac,
        48'h0000040059788,
        48'h000007b0346b0,
        48'h000004005978c,
        48'h000007b0346b4,
        48'h0000040059790,
        48'h000007b0346b8,
        48'h0000040059794,
        48'h000007b0346bc,
        48'h00000400e5418,
        48'h000007b0346cc,
        48'h000007b0346cc,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003231c,
        48'h00000400e64a4,
        48'h000007b034694,
        48'h000007b0337fc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034694,
        48'h00000400e5418,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b03474c,
        48'h000007b034748,
        48'h000007b03474c,
        48'h000007b034748,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045bec,
        48'h00000400321e8,
        48'h000004003231c,
        48'h00000400e649c,
        48'h00000400e64a4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003231c,
        48'h00000400e64bc,
        48'h000007b034690,
        48'h00000400e64bc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b0346c4,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b0346c4,
        48'h000007b03477c,
        48'h000007b034778,
        48'h000007b034754,
        48'h000007b034750,
        48'h000007b0346a8,
        48'h000007b034690,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b03480c,
        48'h000007b034808,
        48'h000007b03480c,
        48'h000007b034808,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045b48,
        48'h00000400321e8,
        48'h0000040032278,
        48'h0000040073cc4,
        48'h0000040073ccc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032278,
        48'h0000040076190,
        48'h000007b034750,
        48'h0000040076190,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0346b8,
        48'h000007b034750,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b03480c,
        48'h000007b034808,
        48'h000007b03480c,
        48'h000007b034808,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045b50,
        48'h00000400321e8,
        48'h0000040032280,
        48'h0000040096fd4,
        48'h0000040096fdc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032280,
        48'h00000400994a0,
        48'h000007b034778,
        48'h00000400994a0,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034534,
        48'h000007b034778,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b034804,
        48'h0000040020544,
        48'h0000040020764,
        48'h0000040020820,
        48'h0000040020544,
        48'h000007b03480c,
        48'h000007b03480c,
        48'h0000040020544,
        48'h000007b03488c,
        48'h000007b03488c,
        48'h000007b034904,
        48'h0000040020054,
        48'h000007b034904,
        48'h0000040020050,
        48'h0000040020014,
        48'h0000040020734,
        48'h0000040020004,
        48'h000004001fffc,
        48'h000004001ffe0,
        48'h000004001fffc,
        48'h000004002000c,
        48'h000004002000c,
        48'h0000040020014,
        48'h0000040020014,
        48'h0000040020018,
        48'h0000040020018,
        48'h000004002001c,
        48'h000004002001c,
        48'h0000040020058,
        48'h0000040020008,
        48'h00000400207e8,
        48'h00000400207bc,
        48'h000007b034804,
        48'h0000040020054,
        48'h000007b0337fc,
        48'h000004002004c,
        48'h000004002004c,
        48'h000004002076c,
        48'h0000040020774,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h00000400207bc,
        48'h0000040020500,
        48'h000004003220c,
        48'h000007b034534,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040020528,
        48'h0000040032250,
        48'h000004003223c,
        48'h000007b034534,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040020528,
        48'h0000040032250,
        48'h0000040032238,
        48'h0000040020528,
        48'h000004002052c,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032250,
        48'h000004003223c,
        48'h000004003223c,
        48'h000004002052c,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032254,
        48'h000004003bea4,
        48'h000004003bea4,
        48'h000004002052c,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032258,
        48'h0000040045b0c,
        48'h0000040045b0c,
        48'h000004002052c,
        48'h0000040020530,
        48'h0000040020530,
        48'h0000040020534,
        48'h0000040020534,
        48'h0000040020500,
        48'h00000400321ec,
        48'h000007b034534,
        48'h000004003bfb4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034804,
        48'h000007b034754,
        48'h000007b034804,
        48'h000007b034804,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000007b034534,
        48'h000004003234c,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h000007b034778,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b034784,
        48'h000007b034780,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b034784,
        48'h000007b034780,
        48'h000007b03483c,
        48'h000007b034754,
        48'h000007b0337fc,
        48'h000007b0346a8,
        48'h000007b034690,
        48'h000007b03484c,
        48'h000007b034848,
        48'h000007b03484c,
        48'h000007b034848,
        48'h000007b0348cc,
        48'h000007b0348c8,
        48'h000007b0348cc,
        48'h000007b0348c8,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045b48,
        48'h00000400321e8,
        48'h0000040032278,
        48'h0000040073cc4,
        48'h0000040073ccc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032278,
        48'h0000040076190,
        48'h000007b03483c,
        48'h0000040076190,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0346b4,
        48'h000007b03483c,
        48'h000007b03484c,
        48'h000007b034848,
        48'h000007b034844,
        48'h000007b03484c,
        48'h000007b034848,
        48'h000007b034844,
        48'h000007b0348cc,
        48'h000007b0348c8,
        48'h000007b0348cc,
        48'h000007b0348c8,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045b4c,
        48'h00000400321e8,
        48'h000004003227c,
        48'h000004007f88c,
        48'h000004007f894,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003227c,
        48'h00000400207bc,
        48'h0000040020784,
        48'h0000040020764,
        48'h0000040020820,
        48'h000007b0337fc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h000007b034834,
        48'h000007b0337fc,
        48'h000007b034698,
        48'h000007b034754,
        48'h000007b034698,
        48'h0000040020464,
        48'h000007b0337fc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034754,
        48'h00000400edc7c,
        48'h00000400edc80,
        48'h000007b034534,
        48'h0000040020468,
        48'h000007b03478c,
        48'h000007b034788,
        48'h000007b03478c,
        48'h000007b034788,
        48'h0000040020500,
        48'h00000400321ec,
        48'h000004003bfb4,
        48'h0000040020500,
        48'h00000400321ec,
        48'h000004003bfb4,
        48'h00000400edc88,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c1c,
        48'h0000040045c1c,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034778,
        48'h000007b0337fc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h00000400e53f8,
        48'h00000400e53f4,
        48'h000007b0337fc,
        48'h00000400e5400,
        48'h000007b034534,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b03473c,
        48'h000007b03474c,
        48'h000007b034748,
        48'h000007b034744,
        48'h000007b03474c,
        48'h000007b034748,
        48'h000007b034744,
        48'h000007b0337fc,
        48'h000007b03473c,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045bf4,
        48'h00000400321e8,
        48'h0000040032324,
        48'h00000400e6aac,
        48'h00000400e6ab4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b03473c,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032324,
        48'h00000400e6acc,
        48'h00000400e6acc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h00000400e5408,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b03473c,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003232c,
        48'h00000400e70c0,
        48'h000007b03474c,
        48'h000007b034748,
        48'h000007b034744,
        48'h000007b03474c,
        48'h000007b034748,
        48'h000007b034744,
        48'h000007b0337fc,
        48'h000007b03473c,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045bfc,
        48'h00000400321e8,
        48'h000004003232c,
        48'h00000400e70bc,
        48'h00000400e70c4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003232c,
        48'h00000400e70d8,
        48'h00000400e70d8,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h00000400e5404,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b03473c,
        48'h000007b03474c,
        48'h000007b034748,
        48'h000007b034744,
        48'h000007b03474c,
        48'h000007b034748,
        48'h000007b034744,
        48'h000007b0337fc,
        48'h000007b03473c,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045bf8,
        48'h00000400321e8,
        48'h0000040032328,
        48'h00000400e6db4,
        48'h00000400e6dbc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b03473c,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032328,
        48'h00000400e6dd4,
        48'h00000400e6dd4,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h00000400597c0,
        48'h00000400e53d4,
        48'h00000400e53c8,
        48'h00000400e5414,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b0346cc,
        48'h000007b0346c8,
        48'h000007b03474c,
        48'h000007b034748,
        48'h000007b03474c,
        48'h000007b034748,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321f0,
        48'h0000040045c08,
        48'h00000400321e8,
        48'h0000040032338,
        48'h00000400ed254,
        48'h00000400ed25c,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h0000040032338,
        48'h00000400ed274,
        48'h000007b03468c,
        48'h00000400ed274,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b03468c,
        48'h000007b034534,
        48'h000007b0346cc,
        48'h000007b0346cc,
        48'h0000040020530,
        48'h0000040020504,
        48'h000007b0337fc,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003234c,
        48'h000007b034688,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034534,
        48'h000007b0346cc,
        48'h000007b0346cc,
        48'h0000040020504,
        48'h0000040020500,
        48'h00000400321e8,
        48'h000004003234c,
        48'h00000400edc84,
        48'h000007b034684,
        48'h000007b0337fc,
        48'h000007b0337fc,
        48'h0000040020760,
        48'h0000040020760,
        48'h000007b034688,
        48'h000007b034684,
        48'h00000400edc98,
        48'h000007b034684,
        48'h00000400edca0,
        48'h000007b034684,
        48'h00000400edca8,
        48'h000007b034684,
        48'h00000400edcb0,
        48'h000007b034684,
        48'h00000400edcb8,
        48'h000007b034684,
        48'h00000400edcc0,
        48'h000007b034684,
        48'h00000400edcc8,
        48'h000007b034684,
        48'h00000400edcd0,
        48'h000007b034684,
        48'h00000400edcd8,
        48'h000007b034684,
        48'h00000400edce0,
        48'h000007b034684,
        48'h00000400edce8,
        48'h000007b034684,
        48'h00000400edcf0,
        48'h000007b034684,
        48'h00000400edcf8,
        48'h000007b034684,
        48'h00000400edd00,
        48'h000007b034684,
        48'h00000400edd08,
        48'h000007b034684,
        48'h00000400edd10,
        48'h000007b034684,
        48'h00000400edd18,
        48'h000007b034684,
        48'h00000400edd20,
        48'h000007b034684,
        48'h00000400edd28,
        48'h000007b034684,
        48'h00000400edd30,
        48'h000007b034684,
        48'h00000400edd38,
        48'h000007b034684,
        48'h00000400edd40,
        48'h000007b034684,
        48'h00000400edd48,
        48'h000007b034684,
        48'h00000400edd50,
        48'h000007b034684,
        48'h00000400edd58,
        48'h000007b034684,
        48'h00000400edd60,
        48'h000007b034684,
        48'h00000400edd68,
        48'h000007b034684,
        48'h00000400edd70,
        48'h000007b034684,
        48'h00000400edd78,
        48'h000007b034684,
        48'h00000400edd80,
        48'h000007b034684,
        48'h00000400edd88,
        48'h000007b034684,
        48'h00000400edd90,
        48'h000007b034684,
        48'h00000400edd98,
        48'h000007b034684,
        48'h00000400edda0,
        48'h000007b034684,
        48'h00000400edda8,
        48'h000007b034684,
        48'h00000400eddb0,
        48'h000007b034684,
        48'h00000400eddb8,
        48'h000007b034684,
        48'h00000400eddc0,
        48'h000007b034684,
        48'h00000400eddc8,
        48'h000007b034684,
        48'h00000400eddd0,
        48'h000007b034684,
        48'h00000400eddd8,
        48'h000007b034684
        };
endmodule
